######################################################################
#  Copyright 1998 - 2023 Dolphin Technology, Inc.                    #
#  This memory compiler and any data created by it are proprietary   #
#  and confidential information of Dolphin Technology, Inc. and      #
#  can only be used or viewed with written permission from           #
#  Dolphin Technology, Inc.                                          #
#  tsmc16nmffcll with hvt, version 1p1p61 Rev_1.5                    #
######################################################################

VERSION 5.4 ;
VERSION 5.5 ;
VERSION 5.6 ;
VERSION 5.7 ;
NAMESCASESENSITIVE ON ;
SITE dti_1pr_ll_tm16ffcllhvt_64x128_1ww2x_m_shc
  CLASS CORE ; 
  SIZE 26.966 by 72.096 ;
  SYMMETRY X Y ; 
END dti_1pr_ll_tm16ffcllhvt_64x128_1ww2x_m_shc
MACRO dti_1pr_ll_tm16ffcllhvt_64x128_1ww2x_m_shc
  CLASS BLOCK ; 
  FOREIGN dti_1pr_ll_tm16ffcllhvt_64x128_1ww2x_m_shc ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.966 by 72.096 ;
  SYMMETRY X Y ; 
  SITE dti_1pr_ll_tm16ffcllhvt_64x128_1ww2x_m_shc ;
  PIN DO[0]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 0.8530 26.9660 0.8910 ;
      LAYER M3 ;
      RECT 26.9020 0.8530 26.9660 0.8910 ;
    END
  END DO[0]
  PIN DI[0]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 0.9230 26.9660 0.9610 ;
      LAYER M3 ;
      RECT 26.9020 0.9230 26.9660 0.9610 ;
    END
  END DI[0]
  PIN DI[1]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 1.0550 26.9660 1.0930 ;
      LAYER M3 ;
      RECT 26.9020 1.0550 26.9660 1.0930 ;
    END
  END DI[1]
  PIN DO[1]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 1.1250 26.9660 1.1630 ;
      LAYER M3 ;
      RECT 26.9020 1.1250 26.9660 1.1630 ;
    END
  END DO[1]
  PIN DO[2]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 1.8130 26.9660 1.8510 ;
      LAYER M3 ;
      RECT 26.9020 1.8130 26.9660 1.8510 ;
    END
  END DO[2]
  PIN DI[2]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 1.8830 26.9660 1.9210 ;
      LAYER M3 ;
      RECT 26.9020 1.8830 26.9660 1.9210 ;
    END
  END DI[2]
  PIN DI[3]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 2.0150 26.9660 2.0530 ;
      LAYER M3 ;
      RECT 26.9020 2.0150 26.9660 2.0530 ;
    END
  END DI[3]
  PIN DO[3]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 2.0850 26.9660 2.1230 ;
      LAYER M3 ;
      RECT 26.9020 2.0850 26.9660 2.1230 ;
    END
  END DO[3]
  PIN DO[4]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 2.7730 26.9660 2.8110 ;
      LAYER M3 ;
      RECT 26.9020 2.7730 26.9660 2.8110 ;
    END
  END DO[4]
  PIN DI[4]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 2.8430 26.9660 2.8810 ;
      LAYER M3 ;
      RECT 26.9020 2.8430 26.9660 2.8810 ;
    END
  END DI[4]
  PIN DI[5]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 2.9750 26.9660 3.0130 ;
      LAYER M3 ;
      RECT 26.9020 2.9750 26.9660 3.0130 ;
    END
  END DI[5]
  PIN DO[5]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 3.0450 26.9660 3.0830 ;
      LAYER M3 ;
      RECT 26.9020 3.0450 26.9660 3.0830 ;
    END
  END DO[5]
  PIN DO[6]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 3.7330 26.9660 3.7710 ;
      LAYER M3 ;
      RECT 26.9020 3.7330 26.9660 3.7710 ;
    END
  END DO[6]
  PIN DI[6]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 3.8030 26.9660 3.8410 ;
      LAYER M3 ;
      RECT 26.9020 3.8030 26.9660 3.8410 ;
    END
  END DI[6]
  PIN DI[7]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 3.9350 26.9660 3.9730 ;
      LAYER M3 ;
      RECT 26.9020 3.9350 26.9660 3.9730 ;
    END
  END DI[7]
  PIN DO[7]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 4.0050 26.9660 4.0430 ;
      LAYER M3 ;
      RECT 26.9020 4.0050 26.9660 4.0430 ;
    END
  END DO[7]
  PIN DO[8]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 4.6930 26.9660 4.7310 ;
      LAYER M3 ;
      RECT 26.9020 4.6930 26.9660 4.7310 ;
    END
  END DO[8]
  PIN DI[8]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 4.7630 26.9660 4.8010 ;
      LAYER M3 ;
      RECT 26.9020 4.7630 26.9660 4.8010 ;
    END
  END DI[8]
  PIN DI[9]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 4.8950 26.9660 4.9330 ;
      LAYER M3 ;
      RECT 26.9020 4.8950 26.9660 4.9330 ;
    END
  END DI[9]
  PIN DO[9]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 4.9650 26.9660 5.0030 ;
      LAYER M3 ;
      RECT 26.9020 4.9650 26.9660 5.0030 ;
    END
  END DO[9]
  PIN DO[10]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 5.6530 26.9660 5.6910 ;
      LAYER M3 ;
      RECT 26.9020 5.6530 26.9660 5.6910 ;
    END
  END DO[10]
  PIN DI[10]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 5.7230 26.9660 5.7610 ;
      LAYER M3 ;
      RECT 26.9020 5.7230 26.9660 5.7610 ;
    END
  END DI[10]
  PIN DI[11]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 5.8550 26.9660 5.8930 ;
      LAYER M3 ;
      RECT 26.9020 5.8550 26.9660 5.8930 ;
    END
  END DI[11]
  PIN DO[11]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 5.9250 26.9660 5.9630 ;
      LAYER M3 ;
      RECT 26.9020 5.9250 26.9660 5.9630 ;
    END
  END DO[11]
  PIN DO[12]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 6.6130 26.9660 6.6510 ;
      LAYER M3 ;
      RECT 26.9020 6.6130 26.9660 6.6510 ;
    END
  END DO[12]
  PIN DI[12]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 6.6830 26.9660 6.7210 ;
      LAYER M3 ;
      RECT 26.9020 6.6830 26.9660 6.7210 ;
    END
  END DI[12]
  PIN DI[13]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 6.8150 26.9660 6.8530 ;
      LAYER M3 ;
      RECT 26.9020 6.8150 26.9660 6.8530 ;
    END
  END DI[13]
  PIN DO[13]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 6.8850 26.9660 6.9230 ;
      LAYER M3 ;
      RECT 26.9020 6.8850 26.9660 6.9230 ;
    END
  END DO[13]
  PIN DO[14]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 7.5730 26.9660 7.6110 ;
      LAYER M3 ;
      RECT 26.9020 7.5730 26.9660 7.6110 ;
    END
  END DO[14]
  PIN DI[14]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 7.6430 26.9660 7.6810 ;
      LAYER M3 ;
      RECT 26.9020 7.6430 26.9660 7.6810 ;
    END
  END DI[14]
  PIN DI[15]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 7.7750 26.9660 7.8130 ;
      LAYER M3 ;
      RECT 26.9020 7.7750 26.9660 7.8130 ;
    END
  END DI[15]
  PIN DO[15]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 7.8450 26.9660 7.8830 ;
      LAYER M3 ;
      RECT 26.9020 7.8450 26.9660 7.8830 ;
    END
  END DO[15]
  PIN DO[16]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 8.5330 26.9660 8.5710 ;
      LAYER M3 ;
      RECT 26.9020 8.5330 26.9660 8.5710 ;
    END
  END DO[16]
  PIN DI[16]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 8.6030 26.9660 8.6410 ;
      LAYER M3 ;
      RECT 26.9020 8.6030 26.9660 8.6410 ;
    END
  END DI[16]
  PIN DI[17]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 8.7350 26.9660 8.7730 ;
      LAYER M3 ;
      RECT 26.9020 8.7350 26.9660 8.7730 ;
    END
  END DI[17]
  PIN DO[17]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 8.8050 26.9660 8.8430 ;
      LAYER M3 ;
      RECT 26.9020 8.8050 26.9660 8.8430 ;
    END
  END DO[17]
  PIN DO[18]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 9.4930 26.9660 9.5310 ;
      LAYER M3 ;
      RECT 26.9020 9.4930 26.9660 9.5310 ;
    END
  END DO[18]
  PIN DI[18]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 9.5630 26.9660 9.6010 ;
      LAYER M3 ;
      RECT 26.9020 9.5630 26.9660 9.6010 ;
    END
  END DI[18]
  PIN DI[19]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 9.6950 26.9660 9.7330 ;
      LAYER M3 ;
      RECT 26.9020 9.6950 26.9660 9.7330 ;
    END
  END DI[19]
  PIN DO[19]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 9.7650 26.9660 9.8030 ;
      LAYER M3 ;
      RECT 26.9020 9.7650 26.9660 9.8030 ;
    END
  END DO[19]
  PIN DO[20]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 10.4530 26.9660 10.4910 ;
      LAYER M3 ;
      RECT 26.9020 10.4530 26.9660 10.4910 ;
    END
  END DO[20]
  PIN DI[20]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 10.5230 26.9660 10.5610 ;
      LAYER M3 ;
      RECT 26.9020 10.5230 26.9660 10.5610 ;
    END
  END DI[20]
  PIN DI[21]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 10.6550 26.9660 10.6930 ;
      LAYER M3 ;
      RECT 26.9020 10.6550 26.9660 10.6930 ;
    END
  END DI[21]
  PIN DO[21]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 10.7250 26.9660 10.7630 ;
      LAYER M3 ;
      RECT 26.9020 10.7250 26.9660 10.7630 ;
    END
  END DO[21]
  PIN DO[22]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 11.4130 26.9660 11.4510 ;
      LAYER M3 ;
      RECT 26.9020 11.4130 26.9660 11.4510 ;
    END
  END DO[22]
  PIN DI[22]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 11.4830 26.9660 11.5210 ;
      LAYER M3 ;
      RECT 26.9020 11.4830 26.9660 11.5210 ;
    END
  END DI[22]
  PIN DI[23]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 11.6150 26.9660 11.6530 ;
      LAYER M3 ;
      RECT 26.9020 11.6150 26.9660 11.6530 ;
    END
  END DI[23]
  PIN DO[23]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 11.6850 26.9660 11.7230 ;
      LAYER M3 ;
      RECT 26.9020 11.6850 26.9660 11.7230 ;
    END
  END DO[23]
  PIN DO[24]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 12.3730 26.9660 12.4110 ;
      LAYER M3 ;
      RECT 26.9020 12.3730 26.9660 12.4110 ;
    END
  END DO[24]
  PIN DI[24]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 12.4430 26.9660 12.4810 ;
      LAYER M3 ;
      RECT 26.9020 12.4430 26.9660 12.4810 ;
    END
  END DI[24]
  PIN DI[25]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 12.5750 26.9660 12.6130 ;
      LAYER M3 ;
      RECT 26.9020 12.5750 26.9660 12.6130 ;
    END
  END DI[25]
  PIN DO[25]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 12.6450 26.9660 12.6830 ;
      LAYER M3 ;
      RECT 26.9020 12.6450 26.9660 12.6830 ;
    END
  END DO[25]
  PIN DO[26]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 13.3330 26.9660 13.3710 ;
      LAYER M3 ;
      RECT 26.9020 13.3330 26.9660 13.3710 ;
    END
  END DO[26]
  PIN DI[26]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 13.4030 26.9660 13.4410 ;
      LAYER M3 ;
      RECT 26.9020 13.4030 26.9660 13.4410 ;
    END
  END DI[26]
  PIN DI[27]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 13.5350 26.9660 13.5730 ;
      LAYER M3 ;
      RECT 26.9020 13.5350 26.9660 13.5730 ;
    END
  END DI[27]
  PIN DO[27]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 13.6050 26.9660 13.6430 ;
      LAYER M3 ;
      RECT 26.9020 13.6050 26.9660 13.6430 ;
    END
  END DO[27]
  PIN DO[28]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 14.2930 26.9660 14.3310 ;
      LAYER M3 ;
      RECT 26.9020 14.2930 26.9660 14.3310 ;
    END
  END DO[28]
  PIN DI[28]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 14.3630 26.9660 14.4010 ;
      LAYER M3 ;
      RECT 26.9020 14.3630 26.9660 14.4010 ;
    END
  END DI[28]
  PIN DI[29]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 14.4950 26.9660 14.5330 ;
      LAYER M3 ;
      RECT 26.9020 14.4950 26.9660 14.5330 ;
    END
  END DI[29]
  PIN DO[29]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 14.5650 26.9660 14.6030 ;
      LAYER M3 ;
      RECT 26.9020 14.5650 26.9660 14.6030 ;
    END
  END DO[29]
  PIN DO[30]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 15.2530 26.9660 15.2910 ;
      LAYER M3 ;
      RECT 26.9020 15.2530 26.9660 15.2910 ;
    END
  END DO[30]
  PIN DI[30]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 15.3230 26.9660 15.3610 ;
      LAYER M3 ;
      RECT 26.9020 15.3230 26.9660 15.3610 ;
    END
  END DI[30]
  PIN DI[31]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 15.4550 26.9660 15.4930 ;
      LAYER M3 ;
      RECT 26.9020 15.4550 26.9660 15.4930 ;
    END
  END DI[31]
  PIN DO[31]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 15.5250 26.9660 15.5630 ;
      LAYER M3 ;
      RECT 26.9020 15.5250 26.9660 15.5630 ;
    END
  END DO[31]
  PIN DO[32]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 16.2130 26.9660 16.2510 ;
      LAYER M3 ;
      RECT 26.9020 16.2130 26.9660 16.2510 ;
    END
  END DO[32]
  PIN DI[32]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 16.2830 26.9660 16.3210 ;
      LAYER M3 ;
      RECT 26.9020 16.2830 26.9660 16.3210 ;
    END
  END DI[32]
  PIN DI[33]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 16.4150 26.9660 16.4530 ;
      LAYER M3 ;
      RECT 26.9020 16.4150 26.9660 16.4530 ;
    END
  END DI[33]
  PIN DO[33]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 16.4850 26.9660 16.5230 ;
      LAYER M3 ;
      RECT 26.9020 16.4850 26.9660 16.5230 ;
    END
  END DO[33]
  PIN DO[34]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 17.1730 26.9660 17.2110 ;
      LAYER M3 ;
      RECT 26.9020 17.1730 26.9660 17.2110 ;
    END
  END DO[34]
  PIN DI[34]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 17.2430 26.9660 17.2810 ;
      LAYER M3 ;
      RECT 26.9020 17.2430 26.9660 17.2810 ;
    END
  END DI[34]
  PIN DI[35]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 17.3750 26.9660 17.4130 ;
      LAYER M3 ;
      RECT 26.9020 17.3750 26.9660 17.4130 ;
    END
  END DI[35]
  PIN DO[35]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 17.4450 26.9660 17.4830 ;
      LAYER M3 ;
      RECT 26.9020 17.4450 26.9660 17.4830 ;
    END
  END DO[35]
  PIN DO[36]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 18.1330 26.9660 18.1710 ;
      LAYER M3 ;
      RECT 26.9020 18.1330 26.9660 18.1710 ;
    END
  END DO[36]
  PIN DI[36]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 18.2030 26.9660 18.2410 ;
      LAYER M3 ;
      RECT 26.9020 18.2030 26.9660 18.2410 ;
    END
  END DI[36]
  PIN DI[37]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 18.3350 26.9660 18.3730 ;
      LAYER M3 ;
      RECT 26.9020 18.3350 26.9660 18.3730 ;
    END
  END DI[37]
  PIN DO[37]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 18.4050 26.9660 18.4430 ;
      LAYER M3 ;
      RECT 26.9020 18.4050 26.9660 18.4430 ;
    END
  END DO[37]
  PIN DO[38]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 19.0930 26.9660 19.1310 ;
      LAYER M3 ;
      RECT 26.9020 19.0930 26.9660 19.1310 ;
    END
  END DO[38]
  PIN DI[38]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 19.1630 26.9660 19.2010 ;
      LAYER M3 ;
      RECT 26.9020 19.1630 26.9660 19.2010 ;
    END
  END DI[38]
  PIN DI[39]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 19.2950 26.9660 19.3330 ;
      LAYER M3 ;
      RECT 26.9020 19.2950 26.9660 19.3330 ;
    END
  END DI[39]
  PIN DO[39]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 19.3650 26.9660 19.4030 ;
      LAYER M3 ;
      RECT 26.9020 19.3650 26.9660 19.4030 ;
    END
  END DO[39]
  PIN DO[40]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 20.0530 26.9660 20.0910 ;
      LAYER M3 ;
      RECT 26.9020 20.0530 26.9660 20.0910 ;
    END
  END DO[40]
  PIN DI[40]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 20.1230 26.9660 20.1610 ;
      LAYER M3 ;
      RECT 26.9020 20.1230 26.9660 20.1610 ;
    END
  END DI[40]
  PIN DI[41]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 20.2550 26.9660 20.2930 ;
      LAYER M3 ;
      RECT 26.9020 20.2550 26.9660 20.2930 ;
    END
  END DI[41]
  PIN DO[41]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 20.3250 26.9660 20.3630 ;
      LAYER M3 ;
      RECT 26.9020 20.3250 26.9660 20.3630 ;
    END
  END DO[41]
  PIN DO[42]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 21.0130 26.9660 21.0510 ;
      LAYER M3 ;
      RECT 26.9020 21.0130 26.9660 21.0510 ;
    END
  END DO[42]
  PIN DI[42]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 21.0830 26.9660 21.1210 ;
      LAYER M3 ;
      RECT 26.9020 21.0830 26.9660 21.1210 ;
    END
  END DI[42]
  PIN DI[43]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 21.2150 26.9660 21.2530 ;
      LAYER M3 ;
      RECT 26.9020 21.2150 26.9660 21.2530 ;
    END
  END DI[43]
  PIN DO[43]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 21.2850 26.9660 21.3230 ;
      LAYER M3 ;
      RECT 26.9020 21.2850 26.9660 21.3230 ;
    END
  END DO[43]
  PIN DO[44]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 21.9730 26.9660 22.0110 ;
      LAYER M3 ;
      RECT 26.9020 21.9730 26.9660 22.0110 ;
    END
  END DO[44]
  PIN DI[44]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 22.0430 26.9660 22.0810 ;
      LAYER M3 ;
      RECT 26.9020 22.0430 26.9660 22.0810 ;
    END
  END DI[44]
  PIN DI[45]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 22.1750 26.9660 22.2130 ;
      LAYER M3 ;
      RECT 26.9020 22.1750 26.9660 22.2130 ;
    END
  END DI[45]
  PIN DO[45]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 22.2450 26.9660 22.2830 ;
      LAYER M3 ;
      RECT 26.9020 22.2450 26.9660 22.2830 ;
    END
  END DO[45]
  PIN DO[46]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 22.9330 26.9660 22.9710 ;
      LAYER M3 ;
      RECT 26.9020 22.9330 26.9660 22.9710 ;
    END
  END DO[46]
  PIN DI[46]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 23.0030 26.9660 23.0410 ;
      LAYER M3 ;
      RECT 26.9020 23.0030 26.9660 23.0410 ;
    END
  END DI[46]
  PIN DI[47]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 23.1350 26.9660 23.1730 ;
      LAYER M3 ;
      RECT 26.9020 23.1350 26.9660 23.1730 ;
    END
  END DI[47]
  PIN DO[47]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 23.2050 26.9660 23.2430 ;
      LAYER M3 ;
      RECT 26.9020 23.2050 26.9660 23.2430 ;
    END
  END DO[47]
  PIN DO[48]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 23.8930 26.9660 23.9310 ;
      LAYER M3 ;
      RECT 26.9020 23.8930 26.9660 23.9310 ;
    END
  END DO[48]
  PIN DI[48]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 23.9630 26.9660 24.0010 ;
      LAYER M3 ;
      RECT 26.9020 23.9630 26.9660 24.0010 ;
    END
  END DI[48]
  PIN DI[49]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 24.0950 26.9660 24.1330 ;
      LAYER M3 ;
      RECT 26.9020 24.0950 26.9660 24.1330 ;
    END
  END DI[49]
  PIN DO[49]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 24.1650 26.9660 24.2030 ;
      LAYER M3 ;
      RECT 26.9020 24.1650 26.9660 24.2030 ;
    END
  END DO[49]
  PIN DO[50]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 24.8530 26.9660 24.8910 ;
      LAYER M3 ;
      RECT 26.9020 24.8530 26.9660 24.8910 ;
    END
  END DO[50]
  PIN DI[50]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 24.9230 26.9660 24.9610 ;
      LAYER M3 ;
      RECT 26.9020 24.9230 26.9660 24.9610 ;
    END
  END DI[50]
  PIN DI[51]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 25.0550 26.9660 25.0930 ;
      LAYER M3 ;
      RECT 26.9020 25.0550 26.9660 25.0930 ;
    END
  END DI[51]
  PIN DO[51]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 25.1250 26.9660 25.1630 ;
      LAYER M3 ;
      RECT 26.9020 25.1250 26.9660 25.1630 ;
    END
  END DO[51]
  PIN DO[52]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 25.8130 26.9660 25.8510 ;
      LAYER M3 ;
      RECT 26.9020 25.8130 26.9660 25.8510 ;
    END
  END DO[52]
  PIN DI[52]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 25.8830 26.9660 25.9210 ;
      LAYER M3 ;
      RECT 26.9020 25.8830 26.9660 25.9210 ;
    END
  END DI[52]
  PIN DI[53]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 26.0150 26.9660 26.0530 ;
      LAYER M3 ;
      RECT 26.9020 26.0150 26.9660 26.0530 ;
    END
  END DI[53]
  PIN DO[53]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 26.0850 26.9660 26.1230 ;
      LAYER M3 ;
      RECT 26.9020 26.0850 26.9660 26.1230 ;
    END
  END DO[53]
  PIN DO[54]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 26.7730 26.9660 26.8110 ;
      LAYER M3 ;
      RECT 26.9020 26.7730 26.9660 26.8110 ;
    END
  END DO[54]
  PIN DI[54]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 26.8430 26.9660 26.8810 ;
      LAYER M3 ;
      RECT 26.9020 26.8430 26.9660 26.8810 ;
    END
  END DI[54]
  PIN DI[55]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 26.9750 26.9660 27.0130 ;
      LAYER M3 ;
      RECT 26.9020 26.9750 26.9660 27.0130 ;
    END
  END DI[55]
  PIN DO[55]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 27.0450 26.9660 27.0830 ;
      LAYER M3 ;
      RECT 26.9020 27.0450 26.9660 27.0830 ;
    END
  END DO[55]
  PIN DO[56]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 27.7330 26.9660 27.7710 ;
      LAYER M3 ;
      RECT 26.9020 27.7330 26.9660 27.7710 ;
    END
  END DO[56]
  PIN DI[56]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 27.8030 26.9660 27.8410 ;
      LAYER M3 ;
      RECT 26.9020 27.8030 26.9660 27.8410 ;
    END
  END DI[56]
  PIN DI[57]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 27.9350 26.9660 27.9730 ;
      LAYER M3 ;
      RECT 26.9020 27.9350 26.9660 27.9730 ;
    END
  END DI[57]
  PIN DO[57]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 28.0050 26.9660 28.0430 ;
      LAYER M3 ;
      RECT 26.9020 28.0050 26.9660 28.0430 ;
    END
  END DO[57]
  PIN DO[58]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 28.6930 26.9660 28.7310 ;
      LAYER M3 ;
      RECT 26.9020 28.6930 26.9660 28.7310 ;
    END
  END DO[58]
  PIN DI[58]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 28.7630 26.9660 28.8010 ;
      LAYER M3 ;
      RECT 26.9020 28.7630 26.9660 28.8010 ;
    END
  END DI[58]
  PIN DI[59]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 28.8950 26.9660 28.9330 ;
      LAYER M3 ;
      RECT 26.9020 28.8950 26.9660 28.9330 ;
    END
  END DI[59]
  PIN DO[59]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 28.9650 26.9660 29.0030 ;
      LAYER M3 ;
      RECT 26.9020 28.9650 26.9660 29.0030 ;
    END
  END DO[59]
  PIN DO[60]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 29.6530 26.9660 29.6910 ;
      LAYER M3 ;
      RECT 26.9020 29.6530 26.9660 29.6910 ;
    END
  END DO[60]
  PIN DI[60]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 29.7230 26.9660 29.7610 ;
      LAYER M3 ;
      RECT 26.9020 29.7230 26.9660 29.7610 ;
    END
  END DI[60]
  PIN DI[61]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 29.8550 26.9660 29.8930 ;
      LAYER M3 ;
      RECT 26.9020 29.8550 26.9660 29.8930 ;
    END
  END DI[61]
  PIN DO[61]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 29.9250 26.9660 29.9630 ;
      LAYER M3 ;
      RECT 26.9020 29.9250 26.9660 29.9630 ;
    END
  END DO[61]
  PIN DO[62]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 30.6130 26.9660 30.6510 ;
      LAYER M3 ;
      RECT 26.9020 30.6130 26.9660 30.6510 ;
    END
  END DO[62]
  PIN DI[62]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 30.6830 26.9660 30.7210 ;
      LAYER M3 ;
      RECT 26.9020 30.6830 26.9660 30.7210 ;
    END
  END DI[62]
  PIN DI[63]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 30.8150 26.9660 30.8530 ;
      LAYER M3 ;
      RECT 26.9020 30.8150 26.9660 30.8530 ;
    END
  END DI[63]
  PIN DO[63]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 30.8850 26.9660 30.9230 ;
      LAYER M3 ;
      RECT 26.9020 30.8850 26.9660 30.9230 ;
    END
  END DO[63]
  PIN A[0]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 26.9020 32.4290 26.9660 32.4670 ;
      LAYER M2 ;
      RECT 26.9020 32.4290 26.9660 32.4670 ;
      LAYER M3 ;
      RECT 26.9020 32.4290 26.9660 32.4670 ;
    END
  END A[0]
  PIN A[1]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 26.9020 33.1010 26.9660 33.1390 ;
      LAYER M2 ;
      RECT 26.9020 33.1010 26.9660 33.1390 ;
      LAYER M3 ;
      RECT 26.9020 33.1010 26.9660 33.1390 ;
    END
  END A[1]
  PIN A[2]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 26.9020 34.5730 26.9660 34.6110 ;
      LAYER M2 ;
      RECT 26.9020 34.5730 26.9660 34.6110 ;
      LAYER M3 ;
      RECT 26.9020 34.5730 26.9660 34.6110 ;
    END
  END A[2]
  PIN CLK
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 26.9020 35.0310 26.9660 35.0690 ;
      LAYER M2 ;
      RECT 26.9020 35.0310 26.9660 35.0690 ;
      LAYER M3 ;
      RECT 26.9020 35.0310 26.9660 35.0690 ;
    END
  END CLK
  PIN GWE_N
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 26.9020 35.4430 26.9660 35.4810 ;
      LAYER M2 ;
      RECT 26.9020 35.4430 26.9660 35.4810 ;
      LAYER M3 ;
      RECT 26.9020 35.4430 26.9660 35.4810 ;
    END
  END GWE_N
  PIN CE_N
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT 26.9020 35.5190 26.9660 35.5570 ;
      LAYER M2 ;
      RECT 26.9020 35.5190 26.9660 35.5570 ;
      LAYER M3 ;
      RECT 26.9020 35.5190 26.9660 35.5570 ;
    END
  END CE_N
  PIN A[4]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 26.9020 37.1550 26.9660 37.1930 ;
      LAYER M2 ;
      RECT 26.9020 37.1550 26.9660 37.1930 ;
      LAYER M3 ;
      RECT 26.9020 37.1550 26.9660 37.1930 ;
    END
  END A[4]
  PIN A[5]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 26.9020 37.2610 26.9660 37.2990 ;
      LAYER M2 ;
      RECT 26.9020 37.2610 26.9660 37.2990 ;
      LAYER M3 ;
      RECT 26.9020 37.2610 26.9660 37.2990 ;
    END
  END A[5]
  PIN LKRB_N
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 26.9020 38.1540 26.9660 38.1920 ;
      LAYER M2 ;
      RECT 26.9020 38.1540 26.9660 38.1920 ;
      LAYER M3 ;
      RECT 26.9020 38.1540 26.9660 38.1920 ;
    END
  END LKRB_N
  PIN T_RWM[1]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 26.9020 38.3460 26.9660 38.3840 ;
      LAYER M2 ;
      RECT 26.9020 38.3460 26.9660 38.3840 ;
      LAYER M3 ;
      RECT 26.9020 38.3460 26.9660 38.3840 ;
    END
  END T_RWM[1]
  PIN T_RWM[0]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 26.9020 38.4790 26.9660 38.5170 ;
      LAYER M2 ;
      RECT 26.9020 38.4790 26.9660 38.5170 ;
      LAYER M3 ;
      RECT 26.9020 38.4790 26.9660 38.5170 ;
    END
  END T_RWM[0]
  PIN LOLEAK_N
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 26.9020 38.6170 26.9660 38.6550 ;
      LAYER M2 ;
      RECT 26.9020 38.6170 26.9660 38.6550 ;
      LAYER M3 ;
      RECT 26.9020 38.6170 26.9660 38.6550 ;
    END
  END LOLEAK_N
  PIN T_RWM[2]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 26.9020 38.9190 26.9660 38.9570 ;
      LAYER M2 ;
      RECT 26.9020 38.9190 26.9660 38.9570 ;
      LAYER M3 ;
      RECT 26.9020 38.9190 26.9660 38.9570 ;
    END
  END T_RWM[2]
  PIN DS[1]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 26.9020 39.0590 26.9660 39.0970 ;
      LAYER M2 ;
      RECT 26.9020 39.0590 26.9660 39.0970 ;
      LAYER M3 ;
      RECT 26.9020 39.0590 26.9660 39.0970 ;
    END
  END DS[1]
  PIN DS[0]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 26.9020 39.1570 26.9660 39.1950 ;
      LAYER M2 ;
      RECT 26.9020 39.1570 26.9660 39.1950 ;
      LAYER M3 ;
      RECT 26.9020 39.1570 26.9660 39.1950 ;
    END
  END DS[0]
  PIN A[3]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 26.9020 39.7840 26.9660 39.8220 ;
      LAYER M2 ;
      RECT 26.9020 39.7840 26.9660 39.8220 ;
      LAYER M3 ;
      RECT 26.9020 39.7840 26.9660 39.8220 ;
    END
  END A[3]
  PIN DO[64]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 41.1730 26.9660 41.2110 ;
      LAYER M3 ;
      RECT 26.9020 41.1730 26.9660 41.2110 ;
    END
  END DO[64]
  PIN DI[64]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 41.2430 26.9660 41.2810 ;
      LAYER M3 ;
      RECT 26.9020 41.2430 26.9660 41.2810 ;
    END
  END DI[64]
  PIN DI[65]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 41.3750 26.9660 41.4130 ;
      LAYER M3 ;
      RECT 26.9020 41.3750 26.9660 41.4130 ;
    END
  END DI[65]
  PIN DO[65]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 41.4450 26.9660 41.4830 ;
      LAYER M3 ;
      RECT 26.9020 41.4450 26.9660 41.4830 ;
    END
  END DO[65]
  PIN DO[66]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 42.1330 26.9660 42.1710 ;
      LAYER M3 ;
      RECT 26.9020 42.1330 26.9660 42.1710 ;
    END
  END DO[66]
  PIN DI[66]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 42.2030 26.9660 42.2410 ;
      LAYER M3 ;
      RECT 26.9020 42.2030 26.9660 42.2410 ;
    END
  END DI[66]
  PIN DI[67]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 42.3350 26.9660 42.3730 ;
      LAYER M3 ;
      RECT 26.9020 42.3350 26.9660 42.3730 ;
    END
  END DI[67]
  PIN DO[67]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 42.4050 26.9660 42.4430 ;
      LAYER M3 ;
      RECT 26.9020 42.4050 26.9660 42.4430 ;
    END
  END DO[67]
  PIN DO[68]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 43.0930 26.9660 43.1310 ;
      LAYER M3 ;
      RECT 26.9020 43.0930 26.9660 43.1310 ;
    END
  END DO[68]
  PIN DI[68]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 43.1630 26.9660 43.2010 ;
      LAYER M3 ;
      RECT 26.9020 43.1630 26.9660 43.2010 ;
    END
  END DI[68]
  PIN DI[69]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 43.2950 26.9660 43.3330 ;
      LAYER M3 ;
      RECT 26.9020 43.2950 26.9660 43.3330 ;
    END
  END DI[69]
  PIN DO[69]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 43.3650 26.9660 43.4030 ;
      LAYER M3 ;
      RECT 26.9020 43.3650 26.9660 43.4030 ;
    END
  END DO[69]
  PIN DO[70]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 44.0530 26.9660 44.0910 ;
      LAYER M3 ;
      RECT 26.9020 44.0530 26.9660 44.0910 ;
    END
  END DO[70]
  PIN DI[70]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 44.1230 26.9660 44.1610 ;
      LAYER M3 ;
      RECT 26.9020 44.1230 26.9660 44.1610 ;
    END
  END DI[70]
  PIN DI[71]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 44.2550 26.9660 44.2930 ;
      LAYER M3 ;
      RECT 26.9020 44.2550 26.9660 44.2930 ;
    END
  END DI[71]
  PIN DO[71]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 44.3250 26.9660 44.3630 ;
      LAYER M3 ;
      RECT 26.9020 44.3250 26.9660 44.3630 ;
    END
  END DO[71]
  PIN DO[72]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 45.0130 26.9660 45.0510 ;
      LAYER M3 ;
      RECT 26.9020 45.0130 26.9660 45.0510 ;
    END
  END DO[72]
  PIN DI[72]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 45.0830 26.9660 45.1210 ;
      LAYER M3 ;
      RECT 26.9020 45.0830 26.9660 45.1210 ;
    END
  END DI[72]
  PIN DI[73]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 45.2150 26.9660 45.2530 ;
      LAYER M3 ;
      RECT 26.9020 45.2150 26.9660 45.2530 ;
    END
  END DI[73]
  PIN DO[73]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 45.2850 26.9660 45.3230 ;
      LAYER M3 ;
      RECT 26.9020 45.2850 26.9660 45.3230 ;
    END
  END DO[73]
  PIN DO[74]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 45.9730 26.9660 46.0110 ;
      LAYER M3 ;
      RECT 26.9020 45.9730 26.9660 46.0110 ;
    END
  END DO[74]
  PIN DI[74]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 46.0430 26.9660 46.0810 ;
      LAYER M3 ;
      RECT 26.9020 46.0430 26.9660 46.0810 ;
    END
  END DI[74]
  PIN DI[75]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 46.1750 26.9660 46.2130 ;
      LAYER M3 ;
      RECT 26.9020 46.1750 26.9660 46.2130 ;
    END
  END DI[75]
  PIN DO[75]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 46.2450 26.9660 46.2830 ;
      LAYER M3 ;
      RECT 26.9020 46.2450 26.9660 46.2830 ;
    END
  END DO[75]
  PIN DO[76]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 46.9330 26.9660 46.9710 ;
      LAYER M3 ;
      RECT 26.9020 46.9330 26.9660 46.9710 ;
    END
  END DO[76]
  PIN DI[76]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 47.0030 26.9660 47.0410 ;
      LAYER M3 ;
      RECT 26.9020 47.0030 26.9660 47.0410 ;
    END
  END DI[76]
  PIN DI[77]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 47.1350 26.9660 47.1730 ;
      LAYER M3 ;
      RECT 26.9020 47.1350 26.9660 47.1730 ;
    END
  END DI[77]
  PIN DO[77]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 47.2050 26.9660 47.2430 ;
      LAYER M3 ;
      RECT 26.9020 47.2050 26.9660 47.2430 ;
    END
  END DO[77]
  PIN DO[78]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 47.8930 26.9660 47.9310 ;
      LAYER M3 ;
      RECT 26.9020 47.8930 26.9660 47.9310 ;
    END
  END DO[78]
  PIN DI[78]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 47.9630 26.9660 48.0010 ;
      LAYER M3 ;
      RECT 26.9020 47.9630 26.9660 48.0010 ;
    END
  END DI[78]
  PIN DI[79]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 48.0950 26.9660 48.1330 ;
      LAYER M3 ;
      RECT 26.9020 48.0950 26.9660 48.1330 ;
    END
  END DI[79]
  PIN DO[79]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 48.1650 26.9660 48.2030 ;
      LAYER M3 ;
      RECT 26.9020 48.1650 26.9660 48.2030 ;
    END
  END DO[79]
  PIN DO[80]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 48.8530 26.9660 48.8910 ;
      LAYER M3 ;
      RECT 26.9020 48.8530 26.9660 48.8910 ;
    END
  END DO[80]
  PIN DI[80]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 48.9230 26.9660 48.9610 ;
      LAYER M3 ;
      RECT 26.9020 48.9230 26.9660 48.9610 ;
    END
  END DI[80]
  PIN DI[81]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 49.0550 26.9660 49.0930 ;
      LAYER M3 ;
      RECT 26.9020 49.0550 26.9660 49.0930 ;
    END
  END DI[81]
  PIN DO[81]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 49.1250 26.9660 49.1630 ;
      LAYER M3 ;
      RECT 26.9020 49.1250 26.9660 49.1630 ;
    END
  END DO[81]
  PIN DO[82]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 49.8130 26.9660 49.8510 ;
      LAYER M3 ;
      RECT 26.9020 49.8130 26.9660 49.8510 ;
    END
  END DO[82]
  PIN DI[82]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 49.8830 26.9660 49.9210 ;
      LAYER M3 ;
      RECT 26.9020 49.8830 26.9660 49.9210 ;
    END
  END DI[82]
  PIN DI[83]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 50.0150 26.9660 50.0530 ;
      LAYER M3 ;
      RECT 26.9020 50.0150 26.9660 50.0530 ;
    END
  END DI[83]
  PIN DO[83]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 50.0850 26.9660 50.1230 ;
      LAYER M3 ;
      RECT 26.9020 50.0850 26.9660 50.1230 ;
    END
  END DO[83]
  PIN DO[84]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 50.7730 26.9660 50.8110 ;
      LAYER M3 ;
      RECT 26.9020 50.7730 26.9660 50.8110 ;
    END
  END DO[84]
  PIN DI[84]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 50.8430 26.9660 50.8810 ;
      LAYER M3 ;
      RECT 26.9020 50.8430 26.9660 50.8810 ;
    END
  END DI[84]
  PIN DI[85]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 50.9750 26.9660 51.0130 ;
      LAYER M3 ;
      RECT 26.9020 50.9750 26.9660 51.0130 ;
    END
  END DI[85]
  PIN DO[85]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 51.0450 26.9660 51.0830 ;
      LAYER M3 ;
      RECT 26.9020 51.0450 26.9660 51.0830 ;
    END
  END DO[85]
  PIN DO[86]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 51.7330 26.9660 51.7710 ;
      LAYER M3 ;
      RECT 26.9020 51.7330 26.9660 51.7710 ;
    END
  END DO[86]
  PIN DI[86]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 51.8030 26.9660 51.8410 ;
      LAYER M3 ;
      RECT 26.9020 51.8030 26.9660 51.8410 ;
    END
  END DI[86]
  PIN DI[87]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 51.9350 26.9660 51.9730 ;
      LAYER M3 ;
      RECT 26.9020 51.9350 26.9660 51.9730 ;
    END
  END DI[87]
  PIN DO[87]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 52.0050 26.9660 52.0430 ;
      LAYER M3 ;
      RECT 26.9020 52.0050 26.9660 52.0430 ;
    END
  END DO[87]
  PIN DO[88]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 52.6930 26.9660 52.7310 ;
      LAYER M3 ;
      RECT 26.9020 52.6930 26.9660 52.7310 ;
    END
  END DO[88]
  PIN DI[88]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 52.7630 26.9660 52.8010 ;
      LAYER M3 ;
      RECT 26.9020 52.7630 26.9660 52.8010 ;
    END
  END DI[88]
  PIN DI[89]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 52.8950 26.9660 52.9330 ;
      LAYER M3 ;
      RECT 26.9020 52.8950 26.9660 52.9330 ;
    END
  END DI[89]
  PIN DO[89]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 52.9650 26.9660 53.0030 ;
      LAYER M3 ;
      RECT 26.9020 52.9650 26.9660 53.0030 ;
    END
  END DO[89]
  PIN DO[90]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 53.6530 26.9660 53.6910 ;
      LAYER M3 ;
      RECT 26.9020 53.6530 26.9660 53.6910 ;
    END
  END DO[90]
  PIN DI[90]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 53.7230 26.9660 53.7610 ;
      LAYER M3 ;
      RECT 26.9020 53.7230 26.9660 53.7610 ;
    END
  END DI[90]
  PIN DI[91]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 53.8550 26.9660 53.8930 ;
      LAYER M3 ;
      RECT 26.9020 53.8550 26.9660 53.8930 ;
    END
  END DI[91]
  PIN DO[91]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 53.9250 26.9660 53.9630 ;
      LAYER M3 ;
      RECT 26.9020 53.9250 26.9660 53.9630 ;
    END
  END DO[91]
  PIN DO[92]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 54.6130 26.9660 54.6510 ;
      LAYER M3 ;
      RECT 26.9020 54.6130 26.9660 54.6510 ;
    END
  END DO[92]
  PIN DI[92]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 54.6830 26.9660 54.7210 ;
      LAYER M3 ;
      RECT 26.9020 54.6830 26.9660 54.7210 ;
    END
  END DI[92]
  PIN DI[93]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 54.8150 26.9660 54.8530 ;
      LAYER M3 ;
      RECT 26.9020 54.8150 26.9660 54.8530 ;
    END
  END DI[93]
  PIN DO[93]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 54.8850 26.9660 54.9230 ;
      LAYER M3 ;
      RECT 26.9020 54.8850 26.9660 54.9230 ;
    END
  END DO[93]
  PIN DO[94]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 55.5730 26.9660 55.6110 ;
      LAYER M3 ;
      RECT 26.9020 55.5730 26.9660 55.6110 ;
    END
  END DO[94]
  PIN DI[94]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 55.6430 26.9660 55.6810 ;
      LAYER M3 ;
      RECT 26.9020 55.6430 26.9660 55.6810 ;
    END
  END DI[94]
  PIN DI[95]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 55.7750 26.9660 55.8130 ;
      LAYER M3 ;
      RECT 26.9020 55.7750 26.9660 55.8130 ;
    END
  END DI[95]
  PIN DO[95]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 55.8450 26.9660 55.8830 ;
      LAYER M3 ;
      RECT 26.9020 55.8450 26.9660 55.8830 ;
    END
  END DO[95]
  PIN DO[96]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 56.5330 26.9660 56.5710 ;
      LAYER M3 ;
      RECT 26.9020 56.5330 26.9660 56.5710 ;
    END
  END DO[96]
  PIN DI[96]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 56.6030 26.9660 56.6410 ;
      LAYER M3 ;
      RECT 26.9020 56.6030 26.9660 56.6410 ;
    END
  END DI[96]
  PIN DI[97]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 56.7350 26.9660 56.7730 ;
      LAYER M3 ;
      RECT 26.9020 56.7350 26.9660 56.7730 ;
    END
  END DI[97]
  PIN DO[97]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 56.8050 26.9660 56.8430 ;
      LAYER M3 ;
      RECT 26.9020 56.8050 26.9660 56.8430 ;
    END
  END DO[97]
  PIN DO[98]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 57.4930 26.9660 57.5310 ;
      LAYER M3 ;
      RECT 26.9020 57.4930 26.9660 57.5310 ;
    END
  END DO[98]
  PIN DI[98]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 57.5630 26.9660 57.6010 ;
      LAYER M3 ;
      RECT 26.9020 57.5630 26.9660 57.6010 ;
    END
  END DI[98]
  PIN DI[99]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 57.6950 26.9660 57.7330 ;
      LAYER M3 ;
      RECT 26.9020 57.6950 26.9660 57.7330 ;
    END
  END DI[99]
  PIN DO[99]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 57.7650 26.9660 57.8030 ;
      LAYER M3 ;
      RECT 26.9020 57.7650 26.9660 57.8030 ;
    END
  END DO[99]
  PIN DO[100]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 58.4530 26.9660 58.4910 ;
      LAYER M3 ;
      RECT 26.9020 58.4530 26.9660 58.4910 ;
    END
  END DO[100]
  PIN DI[100]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 58.5230 26.9660 58.5610 ;
      LAYER M3 ;
      RECT 26.9020 58.5230 26.9660 58.5610 ;
    END
  END DI[100]
  PIN DI[101]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 58.6550 26.9660 58.6930 ;
      LAYER M3 ;
      RECT 26.9020 58.6550 26.9660 58.6930 ;
    END
  END DI[101]
  PIN DO[101]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 58.7250 26.9660 58.7630 ;
      LAYER M3 ;
      RECT 26.9020 58.7250 26.9660 58.7630 ;
    END
  END DO[101]
  PIN DO[102]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 59.4130 26.9660 59.4510 ;
      LAYER M3 ;
      RECT 26.9020 59.4130 26.9660 59.4510 ;
    END
  END DO[102]
  PIN DI[102]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 59.4830 26.9660 59.5210 ;
      LAYER M3 ;
      RECT 26.9020 59.4830 26.9660 59.5210 ;
    END
  END DI[102]
  PIN DI[103]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 59.6150 26.9660 59.6530 ;
      LAYER M3 ;
      RECT 26.9020 59.6150 26.9660 59.6530 ;
    END
  END DI[103]
  PIN DO[103]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 59.6850 26.9660 59.7230 ;
      LAYER M3 ;
      RECT 26.9020 59.6850 26.9660 59.7230 ;
    END
  END DO[103]
  PIN DO[104]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 60.3730 26.9660 60.4110 ;
      LAYER M3 ;
      RECT 26.9020 60.3730 26.9660 60.4110 ;
    END
  END DO[104]
  PIN DI[104]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 60.4430 26.9660 60.4810 ;
      LAYER M3 ;
      RECT 26.9020 60.4430 26.9660 60.4810 ;
    END
  END DI[104]
  PIN DI[105]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 60.5750 26.9660 60.6130 ;
      LAYER M3 ;
      RECT 26.9020 60.5750 26.9660 60.6130 ;
    END
  END DI[105]
  PIN DO[105]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 60.6450 26.9660 60.6830 ;
      LAYER M3 ;
      RECT 26.9020 60.6450 26.9660 60.6830 ;
    END
  END DO[105]
  PIN DO[106]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 61.3330 26.9660 61.3710 ;
      LAYER M3 ;
      RECT 26.9020 61.3330 26.9660 61.3710 ;
    END
  END DO[106]
  PIN DI[106]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 61.4030 26.9660 61.4410 ;
      LAYER M3 ;
      RECT 26.9020 61.4030 26.9660 61.4410 ;
    END
  END DI[106]
  PIN DI[107]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 61.5350 26.9660 61.5730 ;
      LAYER M3 ;
      RECT 26.9020 61.5350 26.9660 61.5730 ;
    END
  END DI[107]
  PIN DO[107]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 61.6050 26.9660 61.6430 ;
      LAYER M3 ;
      RECT 26.9020 61.6050 26.9660 61.6430 ;
    END
  END DO[107]
  PIN DO[108]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 62.2930 26.9660 62.3310 ;
      LAYER M3 ;
      RECT 26.9020 62.2930 26.9660 62.3310 ;
    END
  END DO[108]
  PIN DI[108]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 62.3630 26.9660 62.4010 ;
      LAYER M3 ;
      RECT 26.9020 62.3630 26.9660 62.4010 ;
    END
  END DI[108]
  PIN DI[109]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 62.4950 26.9660 62.5330 ;
      LAYER M3 ;
      RECT 26.9020 62.4950 26.9660 62.5330 ;
    END
  END DI[109]
  PIN DO[109]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 62.5650 26.9660 62.6030 ;
      LAYER M3 ;
      RECT 26.9020 62.5650 26.9660 62.6030 ;
    END
  END DO[109]
  PIN DO[110]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 63.2530 26.9660 63.2910 ;
      LAYER M3 ;
      RECT 26.9020 63.2530 26.9660 63.2910 ;
    END
  END DO[110]
  PIN DI[110]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 63.3230 26.9660 63.3610 ;
      LAYER M3 ;
      RECT 26.9020 63.3230 26.9660 63.3610 ;
    END
  END DI[110]
  PIN DI[111]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 63.4550 26.9660 63.4930 ;
      LAYER M3 ;
      RECT 26.9020 63.4550 26.9660 63.4930 ;
    END
  END DI[111]
  PIN DO[111]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 63.5250 26.9660 63.5630 ;
      LAYER M3 ;
      RECT 26.9020 63.5250 26.9660 63.5630 ;
    END
  END DO[111]
  PIN DO[112]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 64.2130 26.9660 64.2510 ;
      LAYER M3 ;
      RECT 26.9020 64.2130 26.9660 64.2510 ;
    END
  END DO[112]
  PIN DI[112]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 64.2830 26.9660 64.3210 ;
      LAYER M3 ;
      RECT 26.9020 64.2830 26.9660 64.3210 ;
    END
  END DI[112]
  PIN DI[113]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 64.4150 26.9660 64.4530 ;
      LAYER M3 ;
      RECT 26.9020 64.4150 26.9660 64.4530 ;
    END
  END DI[113]
  PIN DO[113]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 64.4850 26.9660 64.5230 ;
      LAYER M3 ;
      RECT 26.9020 64.4850 26.9660 64.5230 ;
    END
  END DO[113]
  PIN DO[114]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 65.1730 26.9660 65.2110 ;
      LAYER M3 ;
      RECT 26.9020 65.1730 26.9660 65.2110 ;
    END
  END DO[114]
  PIN DI[114]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 65.2430 26.9660 65.2810 ;
      LAYER M3 ;
      RECT 26.9020 65.2430 26.9660 65.2810 ;
    END
  END DI[114]
  PIN DI[115]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 65.3750 26.9660 65.4130 ;
      LAYER M3 ;
      RECT 26.9020 65.3750 26.9660 65.4130 ;
    END
  END DI[115]
  PIN DO[115]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 65.4450 26.9660 65.4830 ;
      LAYER M3 ;
      RECT 26.9020 65.4450 26.9660 65.4830 ;
    END
  END DO[115]
  PIN DO[116]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 66.1330 26.9660 66.1710 ;
      LAYER M3 ;
      RECT 26.9020 66.1330 26.9660 66.1710 ;
    END
  END DO[116]
  PIN DI[116]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 66.2030 26.9660 66.2410 ;
      LAYER M3 ;
      RECT 26.9020 66.2030 26.9660 66.2410 ;
    END
  END DI[116]
  PIN DI[117]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 66.3350 26.9660 66.3730 ;
      LAYER M3 ;
      RECT 26.9020 66.3350 26.9660 66.3730 ;
    END
  END DI[117]
  PIN DO[117]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 66.4050 26.9660 66.4430 ;
      LAYER M3 ;
      RECT 26.9020 66.4050 26.9660 66.4430 ;
    END
  END DO[117]
  PIN DO[118]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 67.0930 26.9660 67.1310 ;
      LAYER M3 ;
      RECT 26.9020 67.0930 26.9660 67.1310 ;
    END
  END DO[118]
  PIN DI[118]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 67.1630 26.9660 67.2010 ;
      LAYER M3 ;
      RECT 26.9020 67.1630 26.9660 67.2010 ;
    END
  END DI[118]
  PIN DI[119]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 67.2950 26.9660 67.3330 ;
      LAYER M3 ;
      RECT 26.9020 67.2950 26.9660 67.3330 ;
    END
  END DI[119]
  PIN DO[119]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 67.3650 26.9660 67.4030 ;
      LAYER M3 ;
      RECT 26.9020 67.3650 26.9660 67.4030 ;
    END
  END DO[119]
  PIN DO[120]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 68.0530 26.9660 68.0910 ;
      LAYER M3 ;
      RECT 26.9020 68.0530 26.9660 68.0910 ;
    END
  END DO[120]
  PIN DI[120]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 68.1230 26.9660 68.1610 ;
      LAYER M3 ;
      RECT 26.9020 68.1230 26.9660 68.1610 ;
    END
  END DI[120]
  PIN DI[121]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 68.2550 26.9660 68.2930 ;
      LAYER M3 ;
      RECT 26.9020 68.2550 26.9660 68.2930 ;
    END
  END DI[121]
  PIN DO[121]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 68.3250 26.9660 68.3630 ;
      LAYER M3 ;
      RECT 26.9020 68.3250 26.9660 68.3630 ;
    END
  END DO[121]
  PIN DO[122]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 69.0130 26.9660 69.0510 ;
      LAYER M3 ;
      RECT 26.9020 69.0130 26.9660 69.0510 ;
    END
  END DO[122]
  PIN DI[122]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 69.0830 26.9660 69.1210 ;
      LAYER M3 ;
      RECT 26.9020 69.0830 26.9660 69.1210 ;
    END
  END DI[122]
  PIN DI[123]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 69.2150 26.9660 69.2530 ;
      LAYER M3 ;
      RECT 26.9020 69.2150 26.9660 69.2530 ;
    END
  END DI[123]
  PIN DO[123]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 69.2850 26.9660 69.3230 ;
      LAYER M3 ;
      RECT 26.9020 69.2850 26.9660 69.3230 ;
    END
  END DO[123]
  PIN DO[124]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 69.9730 26.9660 70.0110 ;
      LAYER M3 ;
      RECT 26.9020 69.9730 26.9660 70.0110 ;
    END
  END DO[124]
  PIN DI[124]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 70.0430 26.9660 70.0810 ;
      LAYER M3 ;
      RECT 26.9020 70.0430 26.9660 70.0810 ;
    END
  END DI[124]
  PIN DI[125]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 70.1750 26.9660 70.2130 ;
      LAYER M3 ;
      RECT 26.9020 70.1750 26.9660 70.2130 ;
    END
  END DI[125]
  PIN DO[125]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 70.2450 26.9660 70.2830 ;
      LAYER M3 ;
      RECT 26.9020 70.2450 26.9660 70.2830 ;
    END
  END DO[125]
  PIN DO[126]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 70.9330 26.9660 70.9710 ;
      LAYER M3 ;
      RECT 26.9020 70.9330 26.9660 70.9710 ;
    END
  END DO[126]
  PIN DI[126]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 71.0030 26.9660 71.0410 ;
      LAYER M3 ;
      RECT 26.9020 71.0030 26.9660 71.0410 ;
    END
  END DI[126]
  PIN DI[127]
  USE SIGNAL ;
  DIRECTION INPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 71.1350 26.9660 71.1730 ;
      LAYER M3 ;
      RECT 26.9020 71.1350 26.9660 71.1730 ;
    END
  END DI[127]
  PIN DO[127]
  USE SIGNAL ;
  DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      RECT 26.9020 71.2050 26.9660 71.2430 ;
      LAYER M3 ;
      RECT 26.9020 71.2050 26.9660 71.2430 ;
    END
  END DO[127]
  OBS
    LAYER M1 ;
    RECT 0.5500 0.5500 26.4160 71.5460 ;
    RECT 26.4160 0.0000 26.9660 32.3970 ;
    RECT 26.4160 32.3970 26.9020 32.4990 ;
    RECT 26.4160 32.4990 26.9660 33.0690 ;
    RECT 26.4160 33.0690 26.9020 33.1710 ;
    RECT 26.4160 33.1710 26.9660 34.5410 ;
    RECT 26.4160 34.5410 26.9020 34.6430 ;
    RECT 26.4160 34.6430 26.9660 34.9990 ;
    RECT 26.4160 34.9990 26.9020 35.1010 ;
    RECT 26.4160 35.1010 26.9660 35.4110 ;
    RECT 26.4160 35.4110 26.9020 35.5130 ;
    RECT 26.4160 35.5130 26.9020 35.5890 ;
    RECT 26.4160 35.5890 26.9660 37.1230 ;
    RECT 26.4160 37.1230 26.9020 37.2250 ;
    RECT 26.4160 37.2250 26.9020 37.3310 ;
    RECT 26.4160 37.3310 26.9660 38.1220 ;
    RECT 26.4160 38.1220 26.9020 38.2240 ;
    RECT 26.4160 38.2240 26.9660 38.3140 ;
    RECT 26.4160 38.3140 26.9020 38.4160 ;
    RECT 26.4160 38.4160 26.9020 38.5490 ;
    RECT 26.4160 38.5490 26.9020 38.6870 ;
    RECT 26.4160 38.6870 26.9660 38.8870 ;
    RECT 26.4160 38.8870 26.9020 38.9890 ;
    RECT 26.4160 38.9890 26.9020 39.1290 ;
    RECT 26.4160 39.1290 26.9020 39.2270 ;
    RECT 26.4160 39.2270 26.9660 39.7520 ;
    RECT 26.4160 39.7520 26.9020 39.8540 ;
    RECT 26.4160 39.8540 26.9660 72.0960 ;
    RECT 0.0000 0.0000 0.5500 72.0960 ;
    RECT 0.0000 0.0000 26.9660 0.5500 ;
    RECT 0.0000 71.5460 26.9660 72.0960 ;
    LAYER M2 ;
    RECT 0.5500 0.5500 26.4160 71.5460 ;
    RECT 26.4160 0.0000 26.9660 0.8210 ;
    RECT 26.4160 0.8210 26.9020 0.9230 ;
    RECT 26.4160 0.9230 26.9020 0.9930 ;
    RECT 26.4160 0.9930 26.9020 1.1250 ;
    RECT 26.4160 1.1250 26.9020 1.1950 ;
    RECT 26.4160 1.1950 26.9660 1.7810 ;
    RECT 26.4160 1.7810 26.9020 1.8830 ;
    RECT 26.4160 1.8830 26.9020 1.9530 ;
    RECT 26.4160 1.9530 26.9020 2.0850 ;
    RECT 26.4160 2.0850 26.9020 2.1550 ;
    RECT 26.4160 2.1550 26.9660 2.7410 ;
    RECT 26.4160 2.7410 26.9020 2.8430 ;
    RECT 26.4160 2.8430 26.9020 2.9130 ;
    RECT 26.4160 2.9130 26.9020 3.0450 ;
    RECT 26.4160 3.0450 26.9020 3.1150 ;
    RECT 26.4160 3.1150 26.9660 3.7010 ;
    RECT 26.4160 3.7010 26.9020 3.8030 ;
    RECT 26.4160 3.8030 26.9020 3.8730 ;
    RECT 26.4160 3.8730 26.9020 4.0050 ;
    RECT 26.4160 4.0050 26.9020 4.0750 ;
    RECT 26.4160 4.0750 26.9660 4.6610 ;
    RECT 26.4160 4.6610 26.9020 4.7630 ;
    RECT 26.4160 4.7630 26.9020 4.8330 ;
    RECT 26.4160 4.8330 26.9020 4.9650 ;
    RECT 26.4160 4.9650 26.9020 5.0350 ;
    RECT 26.4160 5.0350 26.9660 5.6210 ;
    RECT 26.4160 5.6210 26.9020 5.7230 ;
    RECT 26.4160 5.7230 26.9020 5.7930 ;
    RECT 26.4160 5.7930 26.9020 5.9250 ;
    RECT 26.4160 5.9250 26.9020 5.9950 ;
    RECT 26.4160 5.9950 26.9660 6.5810 ;
    RECT 26.4160 6.5810 26.9020 6.6830 ;
    RECT 26.4160 6.6830 26.9020 6.7530 ;
    RECT 26.4160 6.7530 26.9020 6.8850 ;
    RECT 26.4160 6.8850 26.9020 6.9550 ;
    RECT 26.4160 6.9550 26.9660 7.5410 ;
    RECT 26.4160 7.5410 26.9020 7.6430 ;
    RECT 26.4160 7.6430 26.9020 7.7130 ;
    RECT 26.4160 7.7130 26.9020 7.8450 ;
    RECT 26.4160 7.8450 26.9020 7.9150 ;
    RECT 26.4160 7.9150 26.9660 8.5010 ;
    RECT 26.4160 8.5010 26.9020 8.6030 ;
    RECT 26.4160 8.6030 26.9020 8.6730 ;
    RECT 26.4160 8.6730 26.9020 8.8050 ;
    RECT 26.4160 8.8050 26.9020 8.8750 ;
    RECT 26.4160 8.8750 26.9660 9.4610 ;
    RECT 26.4160 9.4610 26.9020 9.5630 ;
    RECT 26.4160 9.5630 26.9020 9.6330 ;
    RECT 26.4160 9.6330 26.9020 9.7650 ;
    RECT 26.4160 9.7650 26.9020 9.8350 ;
    RECT 26.4160 9.8350 26.9660 10.4210 ;
    RECT 26.4160 10.4210 26.9020 10.5230 ;
    RECT 26.4160 10.5230 26.9020 10.5930 ;
    RECT 26.4160 10.5930 26.9020 10.7250 ;
    RECT 26.4160 10.7250 26.9020 10.7950 ;
    RECT 26.4160 10.7950 26.9660 11.3810 ;
    RECT 26.4160 11.3810 26.9020 11.4830 ;
    RECT 26.4160 11.4830 26.9020 11.5530 ;
    RECT 26.4160 11.5530 26.9020 11.6850 ;
    RECT 26.4160 11.6850 26.9020 11.7550 ;
    RECT 26.4160 11.7550 26.9660 12.3410 ;
    RECT 26.4160 12.3410 26.9020 12.4430 ;
    RECT 26.4160 12.4430 26.9020 12.5130 ;
    RECT 26.4160 12.5130 26.9020 12.6450 ;
    RECT 26.4160 12.6450 26.9020 12.7150 ;
    RECT 26.4160 12.7150 26.9660 13.3010 ;
    RECT 26.4160 13.3010 26.9020 13.4030 ;
    RECT 26.4160 13.4030 26.9020 13.4730 ;
    RECT 26.4160 13.4730 26.9020 13.6050 ;
    RECT 26.4160 13.6050 26.9020 13.6750 ;
    RECT 26.4160 13.6750 26.9660 14.2610 ;
    RECT 26.4160 14.2610 26.9020 14.3630 ;
    RECT 26.4160 14.3630 26.9020 14.4330 ;
    RECT 26.4160 14.4330 26.9020 14.5650 ;
    RECT 26.4160 14.5650 26.9020 14.6350 ;
    RECT 26.4160 14.6350 26.9660 15.2210 ;
    RECT 26.4160 15.2210 26.9020 15.3230 ;
    RECT 26.4160 15.3230 26.9020 15.3930 ;
    RECT 26.4160 15.3930 26.9020 15.5250 ;
    RECT 26.4160 15.5250 26.9020 15.5950 ;
    RECT 26.4160 15.5950 26.9660 16.1810 ;
    RECT 26.4160 16.1810 26.9020 16.2830 ;
    RECT 26.4160 16.2830 26.9020 16.3530 ;
    RECT 26.4160 16.3530 26.9020 16.4850 ;
    RECT 26.4160 16.4850 26.9020 16.5550 ;
    RECT 26.4160 16.5550 26.9660 17.1410 ;
    RECT 26.4160 17.1410 26.9020 17.2430 ;
    RECT 26.4160 17.2430 26.9020 17.3130 ;
    RECT 26.4160 17.3130 26.9020 17.4450 ;
    RECT 26.4160 17.4450 26.9020 17.5150 ;
    RECT 26.4160 17.5150 26.9660 18.1010 ;
    RECT 26.4160 18.1010 26.9020 18.2030 ;
    RECT 26.4160 18.2030 26.9020 18.2730 ;
    RECT 26.4160 18.2730 26.9020 18.4050 ;
    RECT 26.4160 18.4050 26.9020 18.4750 ;
    RECT 26.4160 18.4750 26.9660 19.0610 ;
    RECT 26.4160 19.0610 26.9020 19.1630 ;
    RECT 26.4160 19.1630 26.9020 19.2330 ;
    RECT 26.4160 19.2330 26.9020 19.3650 ;
    RECT 26.4160 19.3650 26.9020 19.4350 ;
    RECT 26.4160 19.4350 26.9660 20.0210 ;
    RECT 26.4160 20.0210 26.9020 20.1230 ;
    RECT 26.4160 20.1230 26.9020 20.1930 ;
    RECT 26.4160 20.1930 26.9020 20.3250 ;
    RECT 26.4160 20.3250 26.9020 20.3950 ;
    RECT 26.4160 20.3950 26.9660 20.9810 ;
    RECT 26.4160 20.9810 26.9020 21.0830 ;
    RECT 26.4160 21.0830 26.9020 21.1530 ;
    RECT 26.4160 21.1530 26.9020 21.2850 ;
    RECT 26.4160 21.2850 26.9020 21.3550 ;
    RECT 26.4160 21.3550 26.9660 21.9410 ;
    RECT 26.4160 21.9410 26.9020 22.0430 ;
    RECT 26.4160 22.0430 26.9020 22.1130 ;
    RECT 26.4160 22.1130 26.9020 22.2450 ;
    RECT 26.4160 22.2450 26.9020 22.3150 ;
    RECT 26.4160 22.3150 26.9660 22.9010 ;
    RECT 26.4160 22.9010 26.9020 23.0030 ;
    RECT 26.4160 23.0030 26.9020 23.0730 ;
    RECT 26.4160 23.0730 26.9020 23.2050 ;
    RECT 26.4160 23.2050 26.9020 23.2750 ;
    RECT 26.4160 23.2750 26.9660 23.8610 ;
    RECT 26.4160 23.8610 26.9020 23.9630 ;
    RECT 26.4160 23.9630 26.9020 24.0330 ;
    RECT 26.4160 24.0330 26.9020 24.1650 ;
    RECT 26.4160 24.1650 26.9020 24.2350 ;
    RECT 26.4160 24.2350 26.9660 24.8210 ;
    RECT 26.4160 24.8210 26.9020 24.9230 ;
    RECT 26.4160 24.9230 26.9020 24.9930 ;
    RECT 26.4160 24.9930 26.9020 25.1250 ;
    RECT 26.4160 25.1250 26.9020 25.1950 ;
    RECT 26.4160 25.1950 26.9660 25.7810 ;
    RECT 26.4160 25.7810 26.9020 25.8830 ;
    RECT 26.4160 25.8830 26.9020 25.9530 ;
    RECT 26.4160 25.9530 26.9020 26.0850 ;
    RECT 26.4160 26.0850 26.9020 26.1550 ;
    RECT 26.4160 26.1550 26.9660 26.7410 ;
    RECT 26.4160 26.7410 26.9020 26.8430 ;
    RECT 26.4160 26.8430 26.9020 26.9130 ;
    RECT 26.4160 26.9130 26.9020 27.0450 ;
    RECT 26.4160 27.0450 26.9020 27.1150 ;
    RECT 26.4160 27.1150 26.9660 27.7010 ;
    RECT 26.4160 27.7010 26.9020 27.8030 ;
    RECT 26.4160 27.8030 26.9020 27.8730 ;
    RECT 26.4160 27.8730 26.9020 28.0050 ;
    RECT 26.4160 28.0050 26.9020 28.0750 ;
    RECT 26.4160 28.0750 26.9660 28.6610 ;
    RECT 26.4160 28.6610 26.9020 28.7630 ;
    RECT 26.4160 28.7630 26.9020 28.8330 ;
    RECT 26.4160 28.8330 26.9020 28.9650 ;
    RECT 26.4160 28.9650 26.9020 29.0350 ;
    RECT 26.4160 29.0350 26.9660 29.6210 ;
    RECT 26.4160 29.6210 26.9020 29.7230 ;
    RECT 26.4160 29.7230 26.9020 29.7930 ;
    RECT 26.4160 29.7930 26.9020 29.9250 ;
    RECT 26.4160 29.9250 26.9020 29.9950 ;
    RECT 26.4160 29.9950 26.9660 30.5810 ;
    RECT 26.4160 30.5810 26.9020 30.6830 ;
    RECT 26.4160 30.6830 26.9020 30.7530 ;
    RECT 26.4160 30.7530 26.9020 30.8850 ;
    RECT 26.4160 30.8850 26.9020 30.9550 ;
    RECT 26.4160 30.9550 26.9660 32.3970 ;
    RECT 26.4160 32.3970 26.9020 32.4990 ;
    RECT 26.4160 32.4990 26.9660 33.0690 ;
    RECT 26.4160 33.0690 26.9020 33.1710 ;
    RECT 26.4160 33.1710 26.9660 34.5410 ;
    RECT 26.4160 34.5410 26.9020 34.6430 ;
    RECT 26.4160 34.6430 26.9660 34.9990 ;
    RECT 26.4160 34.9990 26.9020 35.1010 ;
    RECT 26.4160 35.1010 26.9660 35.4110 ;
    RECT 26.4160 35.4110 26.9020 35.5130 ;
    RECT 26.4160 35.5130 26.9020 35.5890 ;
    RECT 26.4160 35.5890 26.9660 37.1230 ;
    RECT 26.4160 37.1230 26.9020 37.2250 ;
    RECT 26.4160 37.2250 26.9020 37.3310 ;
    RECT 26.4160 37.3310 26.9660 38.1220 ;
    RECT 26.4160 38.1220 26.9020 38.2240 ;
    RECT 26.4160 38.2240 26.9660 38.3140 ;
    RECT 26.4160 38.3140 26.9020 38.4160 ;
    RECT 26.4160 38.4160 26.9020 38.5490 ;
    RECT 26.4160 38.5490 26.9020 38.6870 ;
    RECT 26.4160 38.6870 26.9660 38.8870 ;
    RECT 26.4160 38.8870 26.9020 38.9890 ;
    RECT 26.4160 38.9890 26.9020 39.1290 ;
    RECT 26.4160 39.1290 26.9020 39.2270 ;
    RECT 26.4160 39.2270 26.9660 39.7520 ;
    RECT 26.4160 39.7520 26.9020 39.8540 ;
    RECT 26.4160 39.8540 26.9660 41.1410 ;
    RECT 26.4160 41.1410 26.9020 41.2430 ;
    RECT 26.4160 41.2430 26.9020 41.3130 ;
    RECT 26.4160 41.3130 26.9020 41.4450 ;
    RECT 26.4160 41.4450 26.9020 41.5150 ;
    RECT 26.4160 41.5150 26.9660 42.1010 ;
    RECT 26.4160 42.1010 26.9020 42.2030 ;
    RECT 26.4160 42.2030 26.9020 42.2730 ;
    RECT 26.4160 42.2730 26.9020 42.4050 ;
    RECT 26.4160 42.4050 26.9020 42.4750 ;
    RECT 26.4160 42.4750 26.9660 43.0610 ;
    RECT 26.4160 43.0610 26.9020 43.1630 ;
    RECT 26.4160 43.1630 26.9020 43.2330 ;
    RECT 26.4160 43.2330 26.9020 43.3650 ;
    RECT 26.4160 43.3650 26.9020 43.4350 ;
    RECT 26.4160 43.4350 26.9660 44.0210 ;
    RECT 26.4160 44.0210 26.9020 44.1230 ;
    RECT 26.4160 44.1230 26.9020 44.1930 ;
    RECT 26.4160 44.1930 26.9020 44.3250 ;
    RECT 26.4160 44.3250 26.9020 44.3950 ;
    RECT 26.4160 44.3950 26.9660 44.9810 ;
    RECT 26.4160 44.9810 26.9020 45.0830 ;
    RECT 26.4160 45.0830 26.9020 45.1530 ;
    RECT 26.4160 45.1530 26.9020 45.2850 ;
    RECT 26.4160 45.2850 26.9020 45.3550 ;
    RECT 26.4160 45.3550 26.9660 45.9410 ;
    RECT 26.4160 45.9410 26.9020 46.0430 ;
    RECT 26.4160 46.0430 26.9020 46.1130 ;
    RECT 26.4160 46.1130 26.9020 46.2450 ;
    RECT 26.4160 46.2450 26.9020 46.3150 ;
    RECT 26.4160 46.3150 26.9660 46.9010 ;
    RECT 26.4160 46.9010 26.9020 47.0030 ;
    RECT 26.4160 47.0030 26.9020 47.0730 ;
    RECT 26.4160 47.0730 26.9020 47.2050 ;
    RECT 26.4160 47.2050 26.9020 47.2750 ;
    RECT 26.4160 47.2750 26.9660 47.8610 ;
    RECT 26.4160 47.8610 26.9020 47.9630 ;
    RECT 26.4160 47.9630 26.9020 48.0330 ;
    RECT 26.4160 48.0330 26.9020 48.1650 ;
    RECT 26.4160 48.1650 26.9020 48.2350 ;
    RECT 26.4160 48.2350 26.9660 48.8210 ;
    RECT 26.4160 48.8210 26.9020 48.9230 ;
    RECT 26.4160 48.9230 26.9020 48.9930 ;
    RECT 26.4160 48.9930 26.9020 49.1250 ;
    RECT 26.4160 49.1250 26.9020 49.1950 ;
    RECT 26.4160 49.1950 26.9660 49.7810 ;
    RECT 26.4160 49.7810 26.9020 49.8830 ;
    RECT 26.4160 49.8830 26.9020 49.9530 ;
    RECT 26.4160 49.9530 26.9020 50.0850 ;
    RECT 26.4160 50.0850 26.9020 50.1550 ;
    RECT 26.4160 50.1550 26.9660 50.7410 ;
    RECT 26.4160 50.7410 26.9020 50.8430 ;
    RECT 26.4160 50.8430 26.9020 50.9130 ;
    RECT 26.4160 50.9130 26.9020 51.0450 ;
    RECT 26.4160 51.0450 26.9020 51.1150 ;
    RECT 26.4160 51.1150 26.9660 51.7010 ;
    RECT 26.4160 51.7010 26.9020 51.8030 ;
    RECT 26.4160 51.8030 26.9020 51.8730 ;
    RECT 26.4160 51.8730 26.9020 52.0050 ;
    RECT 26.4160 52.0050 26.9020 52.0750 ;
    RECT 26.4160 52.0750 26.9660 52.6610 ;
    RECT 26.4160 52.6610 26.9020 52.7630 ;
    RECT 26.4160 52.7630 26.9020 52.8330 ;
    RECT 26.4160 52.8330 26.9020 52.9650 ;
    RECT 26.4160 52.9650 26.9020 53.0350 ;
    RECT 26.4160 53.0350 26.9660 53.6210 ;
    RECT 26.4160 53.6210 26.9020 53.7230 ;
    RECT 26.4160 53.7230 26.9020 53.7930 ;
    RECT 26.4160 53.7930 26.9020 53.9250 ;
    RECT 26.4160 53.9250 26.9020 53.9950 ;
    RECT 26.4160 53.9950 26.9660 54.5810 ;
    RECT 26.4160 54.5810 26.9020 54.6830 ;
    RECT 26.4160 54.6830 26.9020 54.7530 ;
    RECT 26.4160 54.7530 26.9020 54.8850 ;
    RECT 26.4160 54.8850 26.9020 54.9550 ;
    RECT 26.4160 54.9550 26.9660 55.5410 ;
    RECT 26.4160 55.5410 26.9020 55.6430 ;
    RECT 26.4160 55.6430 26.9020 55.7130 ;
    RECT 26.4160 55.7130 26.9020 55.8450 ;
    RECT 26.4160 55.8450 26.9020 55.9150 ;
    RECT 26.4160 55.9150 26.9660 56.5010 ;
    RECT 26.4160 56.5010 26.9020 56.6030 ;
    RECT 26.4160 56.6030 26.9020 56.6730 ;
    RECT 26.4160 56.6730 26.9020 56.8050 ;
    RECT 26.4160 56.8050 26.9020 56.8750 ;
    RECT 26.4160 56.8750 26.9660 57.4610 ;
    RECT 26.4160 57.4610 26.9020 57.5630 ;
    RECT 26.4160 57.5630 26.9020 57.6330 ;
    RECT 26.4160 57.6330 26.9020 57.7650 ;
    RECT 26.4160 57.7650 26.9020 57.8350 ;
    RECT 26.4160 57.8350 26.9660 58.4210 ;
    RECT 26.4160 58.4210 26.9020 58.5230 ;
    RECT 26.4160 58.5230 26.9020 58.5930 ;
    RECT 26.4160 58.5930 26.9020 58.7250 ;
    RECT 26.4160 58.7250 26.9020 58.7950 ;
    RECT 26.4160 58.7950 26.9660 59.3810 ;
    RECT 26.4160 59.3810 26.9020 59.4830 ;
    RECT 26.4160 59.4830 26.9020 59.5530 ;
    RECT 26.4160 59.5530 26.9020 59.6850 ;
    RECT 26.4160 59.6850 26.9020 59.7550 ;
    RECT 26.4160 59.7550 26.9660 60.3410 ;
    RECT 26.4160 60.3410 26.9020 60.4430 ;
    RECT 26.4160 60.4430 26.9020 60.5130 ;
    RECT 26.4160 60.5130 26.9020 60.6450 ;
    RECT 26.4160 60.6450 26.9020 60.7150 ;
    RECT 26.4160 60.7150 26.9660 61.3010 ;
    RECT 26.4160 61.3010 26.9020 61.4030 ;
    RECT 26.4160 61.4030 26.9020 61.4730 ;
    RECT 26.4160 61.4730 26.9020 61.6050 ;
    RECT 26.4160 61.6050 26.9020 61.6750 ;
    RECT 26.4160 61.6750 26.9660 62.2610 ;
    RECT 26.4160 62.2610 26.9020 62.3630 ;
    RECT 26.4160 62.3630 26.9020 62.4330 ;
    RECT 26.4160 62.4330 26.9020 62.5650 ;
    RECT 26.4160 62.5650 26.9020 62.6350 ;
    RECT 26.4160 62.6350 26.9660 63.2210 ;
    RECT 26.4160 63.2210 26.9020 63.3230 ;
    RECT 26.4160 63.3230 26.9020 63.3930 ;
    RECT 26.4160 63.3930 26.9020 63.5250 ;
    RECT 26.4160 63.5250 26.9020 63.5950 ;
    RECT 26.4160 63.5950 26.9660 64.1810 ;
    RECT 26.4160 64.1810 26.9020 64.2830 ;
    RECT 26.4160 64.2830 26.9020 64.3530 ;
    RECT 26.4160 64.3530 26.9020 64.4850 ;
    RECT 26.4160 64.4850 26.9020 64.5550 ;
    RECT 26.4160 64.5550 26.9660 65.1410 ;
    RECT 26.4160 65.1410 26.9020 65.2430 ;
    RECT 26.4160 65.2430 26.9020 65.3130 ;
    RECT 26.4160 65.3130 26.9020 65.4450 ;
    RECT 26.4160 65.4450 26.9020 65.5150 ;
    RECT 26.4160 65.5150 26.9660 66.1010 ;
    RECT 26.4160 66.1010 26.9020 66.2030 ;
    RECT 26.4160 66.2030 26.9020 66.2730 ;
    RECT 26.4160 66.2730 26.9020 66.4050 ;
    RECT 26.4160 66.4050 26.9020 66.4750 ;
    RECT 26.4160 66.4750 26.9660 67.0610 ;
    RECT 26.4160 67.0610 26.9020 67.1630 ;
    RECT 26.4160 67.1630 26.9020 67.2330 ;
    RECT 26.4160 67.2330 26.9020 67.3650 ;
    RECT 26.4160 67.3650 26.9020 67.4350 ;
    RECT 26.4160 67.4350 26.9660 68.0210 ;
    RECT 26.4160 68.0210 26.9020 68.1230 ;
    RECT 26.4160 68.1230 26.9020 68.1930 ;
    RECT 26.4160 68.1930 26.9020 68.3250 ;
    RECT 26.4160 68.3250 26.9020 68.3950 ;
    RECT 26.4160 68.3950 26.9660 68.9810 ;
    RECT 26.4160 68.9810 26.9020 69.0830 ;
    RECT 26.4160 69.0830 26.9020 69.1530 ;
    RECT 26.4160 69.1530 26.9020 69.2850 ;
    RECT 26.4160 69.2850 26.9020 69.3550 ;
    RECT 26.4160 69.3550 26.9660 69.9410 ;
    RECT 26.4160 69.9410 26.9020 70.0430 ;
    RECT 26.4160 70.0430 26.9020 70.1130 ;
    RECT 26.4160 70.1130 26.9020 70.2450 ;
    RECT 26.4160 70.2450 26.9020 70.3150 ;
    RECT 26.4160 70.3150 26.9660 70.9010 ;
    RECT 26.4160 70.9010 26.9020 71.0030 ;
    RECT 26.4160 71.0030 26.9020 71.0730 ;
    RECT 26.4160 71.0730 26.9020 71.2050 ;
    RECT 26.4160 71.2050 26.9020 71.2750 ;
    RECT 26.4160 71.2750 26.9660 72.0960 ;
    RECT 0.0000 0.0000 0.5500 72.0960 ;
    RECT 0.0000 0.0000 26.9660 0.5500 ;
    RECT 0.0000 71.5460 26.9660 72.0960 ;
    LAYER M3 ;
    RECT 0.5500 0.5500 26.4160 71.5460 ;
    RECT 26.4160 0.0000 26.9660 0.8210 ;
    RECT 26.4160 0.8210 26.9020 0.9230 ;
    RECT 26.4160 0.9230 26.9020 0.9930 ;
    RECT 26.4160 0.9930 26.9020 1.1250 ;
    RECT 26.4160 1.1250 26.9020 1.1950 ;
    RECT 26.4160 1.1950 26.9660 1.7810 ;
    RECT 26.4160 1.7810 26.9020 1.8830 ;
    RECT 26.4160 1.8830 26.9020 1.9530 ;
    RECT 26.4160 1.9530 26.9020 2.0850 ;
    RECT 26.4160 2.0850 26.9020 2.1550 ;
    RECT 26.4160 2.1550 26.9660 2.7410 ;
    RECT 26.4160 2.7410 26.9020 2.8430 ;
    RECT 26.4160 2.8430 26.9020 2.9130 ;
    RECT 26.4160 2.9130 26.9020 3.0450 ;
    RECT 26.4160 3.0450 26.9020 3.1150 ;
    RECT 26.4160 3.1150 26.9660 3.7010 ;
    RECT 26.4160 3.7010 26.9020 3.8030 ;
    RECT 26.4160 3.8030 26.9020 3.8730 ;
    RECT 26.4160 3.8730 26.9020 4.0050 ;
    RECT 26.4160 4.0050 26.9020 4.0750 ;
    RECT 26.4160 4.0750 26.9660 4.6610 ;
    RECT 26.4160 4.6610 26.9020 4.7630 ;
    RECT 26.4160 4.7630 26.9020 4.8330 ;
    RECT 26.4160 4.8330 26.9020 4.9650 ;
    RECT 26.4160 4.9650 26.9020 5.0350 ;
    RECT 26.4160 5.0350 26.9660 5.6210 ;
    RECT 26.4160 5.6210 26.9020 5.7230 ;
    RECT 26.4160 5.7230 26.9020 5.7930 ;
    RECT 26.4160 5.7930 26.9020 5.9250 ;
    RECT 26.4160 5.9250 26.9020 5.9950 ;
    RECT 26.4160 5.9950 26.9660 6.5810 ;
    RECT 26.4160 6.5810 26.9020 6.6830 ;
    RECT 26.4160 6.6830 26.9020 6.7530 ;
    RECT 26.4160 6.7530 26.9020 6.8850 ;
    RECT 26.4160 6.8850 26.9020 6.9550 ;
    RECT 26.4160 6.9550 26.9660 7.5410 ;
    RECT 26.4160 7.5410 26.9020 7.6430 ;
    RECT 26.4160 7.6430 26.9020 7.7130 ;
    RECT 26.4160 7.7130 26.9020 7.8450 ;
    RECT 26.4160 7.8450 26.9020 7.9150 ;
    RECT 26.4160 7.9150 26.9660 8.5010 ;
    RECT 26.4160 8.5010 26.9020 8.6030 ;
    RECT 26.4160 8.6030 26.9020 8.6730 ;
    RECT 26.4160 8.6730 26.9020 8.8050 ;
    RECT 26.4160 8.8050 26.9020 8.8750 ;
    RECT 26.4160 8.8750 26.9660 9.4610 ;
    RECT 26.4160 9.4610 26.9020 9.5630 ;
    RECT 26.4160 9.5630 26.9020 9.6330 ;
    RECT 26.4160 9.6330 26.9020 9.7650 ;
    RECT 26.4160 9.7650 26.9020 9.8350 ;
    RECT 26.4160 9.8350 26.9660 10.4210 ;
    RECT 26.4160 10.4210 26.9020 10.5230 ;
    RECT 26.4160 10.5230 26.9020 10.5930 ;
    RECT 26.4160 10.5930 26.9020 10.7250 ;
    RECT 26.4160 10.7250 26.9020 10.7950 ;
    RECT 26.4160 10.7950 26.9660 11.3810 ;
    RECT 26.4160 11.3810 26.9020 11.4830 ;
    RECT 26.4160 11.4830 26.9020 11.5530 ;
    RECT 26.4160 11.5530 26.9020 11.6850 ;
    RECT 26.4160 11.6850 26.9020 11.7550 ;
    RECT 26.4160 11.7550 26.9660 12.3410 ;
    RECT 26.4160 12.3410 26.9020 12.4430 ;
    RECT 26.4160 12.4430 26.9020 12.5130 ;
    RECT 26.4160 12.5130 26.9020 12.6450 ;
    RECT 26.4160 12.6450 26.9020 12.7150 ;
    RECT 26.4160 12.7150 26.9660 13.3010 ;
    RECT 26.4160 13.3010 26.9020 13.4030 ;
    RECT 26.4160 13.4030 26.9020 13.4730 ;
    RECT 26.4160 13.4730 26.9020 13.6050 ;
    RECT 26.4160 13.6050 26.9020 13.6750 ;
    RECT 26.4160 13.6750 26.9660 14.2610 ;
    RECT 26.4160 14.2610 26.9020 14.3630 ;
    RECT 26.4160 14.3630 26.9020 14.4330 ;
    RECT 26.4160 14.4330 26.9020 14.5650 ;
    RECT 26.4160 14.5650 26.9020 14.6350 ;
    RECT 26.4160 14.6350 26.9660 15.2210 ;
    RECT 26.4160 15.2210 26.9020 15.3230 ;
    RECT 26.4160 15.3230 26.9020 15.3930 ;
    RECT 26.4160 15.3930 26.9020 15.5250 ;
    RECT 26.4160 15.5250 26.9020 15.5950 ;
    RECT 26.4160 15.5950 26.9660 16.1810 ;
    RECT 26.4160 16.1810 26.9020 16.2830 ;
    RECT 26.4160 16.2830 26.9020 16.3530 ;
    RECT 26.4160 16.3530 26.9020 16.4850 ;
    RECT 26.4160 16.4850 26.9020 16.5550 ;
    RECT 26.4160 16.5550 26.9660 17.1410 ;
    RECT 26.4160 17.1410 26.9020 17.2430 ;
    RECT 26.4160 17.2430 26.9020 17.3130 ;
    RECT 26.4160 17.3130 26.9020 17.4450 ;
    RECT 26.4160 17.4450 26.9020 17.5150 ;
    RECT 26.4160 17.5150 26.9660 18.1010 ;
    RECT 26.4160 18.1010 26.9020 18.2030 ;
    RECT 26.4160 18.2030 26.9020 18.2730 ;
    RECT 26.4160 18.2730 26.9020 18.4050 ;
    RECT 26.4160 18.4050 26.9020 18.4750 ;
    RECT 26.4160 18.4750 26.9660 19.0610 ;
    RECT 26.4160 19.0610 26.9020 19.1630 ;
    RECT 26.4160 19.1630 26.9020 19.2330 ;
    RECT 26.4160 19.2330 26.9020 19.3650 ;
    RECT 26.4160 19.3650 26.9020 19.4350 ;
    RECT 26.4160 19.4350 26.9660 20.0210 ;
    RECT 26.4160 20.0210 26.9020 20.1230 ;
    RECT 26.4160 20.1230 26.9020 20.1930 ;
    RECT 26.4160 20.1930 26.9020 20.3250 ;
    RECT 26.4160 20.3250 26.9020 20.3950 ;
    RECT 26.4160 20.3950 26.9660 20.9810 ;
    RECT 26.4160 20.9810 26.9020 21.0830 ;
    RECT 26.4160 21.0830 26.9020 21.1530 ;
    RECT 26.4160 21.1530 26.9020 21.2850 ;
    RECT 26.4160 21.2850 26.9020 21.3550 ;
    RECT 26.4160 21.3550 26.9660 21.9410 ;
    RECT 26.4160 21.9410 26.9020 22.0430 ;
    RECT 26.4160 22.0430 26.9020 22.1130 ;
    RECT 26.4160 22.1130 26.9020 22.2450 ;
    RECT 26.4160 22.2450 26.9020 22.3150 ;
    RECT 26.4160 22.3150 26.9660 22.9010 ;
    RECT 26.4160 22.9010 26.9020 23.0030 ;
    RECT 26.4160 23.0030 26.9020 23.0730 ;
    RECT 26.4160 23.0730 26.9020 23.2050 ;
    RECT 26.4160 23.2050 26.9020 23.2750 ;
    RECT 26.4160 23.2750 26.9660 23.8610 ;
    RECT 26.4160 23.8610 26.9020 23.9630 ;
    RECT 26.4160 23.9630 26.9020 24.0330 ;
    RECT 26.4160 24.0330 26.9020 24.1650 ;
    RECT 26.4160 24.1650 26.9020 24.2350 ;
    RECT 26.4160 24.2350 26.9660 24.8210 ;
    RECT 26.4160 24.8210 26.9020 24.9230 ;
    RECT 26.4160 24.9230 26.9020 24.9930 ;
    RECT 26.4160 24.9930 26.9020 25.1250 ;
    RECT 26.4160 25.1250 26.9020 25.1950 ;
    RECT 26.4160 25.1950 26.9660 25.7810 ;
    RECT 26.4160 25.7810 26.9020 25.8830 ;
    RECT 26.4160 25.8830 26.9020 25.9530 ;
    RECT 26.4160 25.9530 26.9020 26.0850 ;
    RECT 26.4160 26.0850 26.9020 26.1550 ;
    RECT 26.4160 26.1550 26.9660 26.7410 ;
    RECT 26.4160 26.7410 26.9020 26.8430 ;
    RECT 26.4160 26.8430 26.9020 26.9130 ;
    RECT 26.4160 26.9130 26.9020 27.0450 ;
    RECT 26.4160 27.0450 26.9020 27.1150 ;
    RECT 26.4160 27.1150 26.9660 27.7010 ;
    RECT 26.4160 27.7010 26.9020 27.8030 ;
    RECT 26.4160 27.8030 26.9020 27.8730 ;
    RECT 26.4160 27.8730 26.9020 28.0050 ;
    RECT 26.4160 28.0050 26.9020 28.0750 ;
    RECT 26.4160 28.0750 26.9660 28.6610 ;
    RECT 26.4160 28.6610 26.9020 28.7630 ;
    RECT 26.4160 28.7630 26.9020 28.8330 ;
    RECT 26.4160 28.8330 26.9020 28.9650 ;
    RECT 26.4160 28.9650 26.9020 29.0350 ;
    RECT 26.4160 29.0350 26.9660 29.6210 ;
    RECT 26.4160 29.6210 26.9020 29.7230 ;
    RECT 26.4160 29.7230 26.9020 29.7930 ;
    RECT 26.4160 29.7930 26.9020 29.9250 ;
    RECT 26.4160 29.9250 26.9020 29.9950 ;
    RECT 26.4160 29.9950 26.9660 30.5810 ;
    RECT 26.4160 30.5810 26.9020 30.6830 ;
    RECT 26.4160 30.6830 26.9020 30.7530 ;
    RECT 26.4160 30.7530 26.9020 30.8850 ;
    RECT 26.4160 30.8850 26.9020 30.9550 ;
    RECT 26.4160 30.9550 26.9660 32.3970 ;
    RECT 26.4160 32.3970 26.9020 32.4990 ;
    RECT 26.4160 32.4990 26.9660 33.0690 ;
    RECT 26.4160 33.0690 26.9020 33.1710 ;
    RECT 26.4160 33.1710 26.9660 34.5410 ;
    RECT 26.4160 34.5410 26.9020 34.6430 ;
    RECT 26.4160 34.6430 26.9660 34.9990 ;
    RECT 26.4160 34.9990 26.9020 35.1010 ;
    RECT 26.4160 35.1010 26.9660 35.4110 ;
    RECT 26.4160 35.4110 26.9020 35.5130 ;
    RECT 26.4160 35.5130 26.9020 35.5890 ;
    RECT 26.4160 35.5890 26.9660 37.1230 ;
    RECT 26.4160 37.1230 26.9020 37.2250 ;
    RECT 26.4160 37.2250 26.9020 37.3310 ;
    RECT 26.4160 37.3310 26.9660 38.1220 ;
    RECT 26.4160 38.1220 26.9020 38.2240 ;
    RECT 26.4160 38.2240 26.9660 38.3140 ;
    RECT 26.4160 38.3140 26.9020 38.4160 ;
    RECT 26.4160 38.4160 26.9020 38.5490 ;
    RECT 26.4160 38.5490 26.9020 38.6870 ;
    RECT 26.4160 38.6870 26.9660 38.8870 ;
    RECT 26.4160 38.8870 26.9020 38.9890 ;
    RECT 26.4160 38.9890 26.9020 39.1290 ;
    RECT 26.4160 39.1290 26.9020 39.2270 ;
    RECT 26.4160 39.2270 26.9660 39.7520 ;
    RECT 26.4160 39.7520 26.9020 39.8540 ;
    RECT 26.4160 39.8540 26.9660 41.1410 ;
    RECT 26.4160 41.1410 26.9020 41.2430 ;
    RECT 26.4160 41.2430 26.9020 41.3130 ;
    RECT 26.4160 41.3130 26.9020 41.4450 ;
    RECT 26.4160 41.4450 26.9020 41.5150 ;
    RECT 26.4160 41.5150 26.9660 42.1010 ;
    RECT 26.4160 42.1010 26.9020 42.2030 ;
    RECT 26.4160 42.2030 26.9020 42.2730 ;
    RECT 26.4160 42.2730 26.9020 42.4050 ;
    RECT 26.4160 42.4050 26.9020 42.4750 ;
    RECT 26.4160 42.4750 26.9660 43.0610 ;
    RECT 26.4160 43.0610 26.9020 43.1630 ;
    RECT 26.4160 43.1630 26.9020 43.2330 ;
    RECT 26.4160 43.2330 26.9020 43.3650 ;
    RECT 26.4160 43.3650 26.9020 43.4350 ;
    RECT 26.4160 43.4350 26.9660 44.0210 ;
    RECT 26.4160 44.0210 26.9020 44.1230 ;
    RECT 26.4160 44.1230 26.9020 44.1930 ;
    RECT 26.4160 44.1930 26.9020 44.3250 ;
    RECT 26.4160 44.3250 26.9020 44.3950 ;
    RECT 26.4160 44.3950 26.9660 44.9810 ;
    RECT 26.4160 44.9810 26.9020 45.0830 ;
    RECT 26.4160 45.0830 26.9020 45.1530 ;
    RECT 26.4160 45.1530 26.9020 45.2850 ;
    RECT 26.4160 45.2850 26.9020 45.3550 ;
    RECT 26.4160 45.3550 26.9660 45.9410 ;
    RECT 26.4160 45.9410 26.9020 46.0430 ;
    RECT 26.4160 46.0430 26.9020 46.1130 ;
    RECT 26.4160 46.1130 26.9020 46.2450 ;
    RECT 26.4160 46.2450 26.9020 46.3150 ;
    RECT 26.4160 46.3150 26.9660 46.9010 ;
    RECT 26.4160 46.9010 26.9020 47.0030 ;
    RECT 26.4160 47.0030 26.9020 47.0730 ;
    RECT 26.4160 47.0730 26.9020 47.2050 ;
    RECT 26.4160 47.2050 26.9020 47.2750 ;
    RECT 26.4160 47.2750 26.9660 47.8610 ;
    RECT 26.4160 47.8610 26.9020 47.9630 ;
    RECT 26.4160 47.9630 26.9020 48.0330 ;
    RECT 26.4160 48.0330 26.9020 48.1650 ;
    RECT 26.4160 48.1650 26.9020 48.2350 ;
    RECT 26.4160 48.2350 26.9660 48.8210 ;
    RECT 26.4160 48.8210 26.9020 48.9230 ;
    RECT 26.4160 48.9230 26.9020 48.9930 ;
    RECT 26.4160 48.9930 26.9020 49.1250 ;
    RECT 26.4160 49.1250 26.9020 49.1950 ;
    RECT 26.4160 49.1950 26.9660 49.7810 ;
    RECT 26.4160 49.7810 26.9020 49.8830 ;
    RECT 26.4160 49.8830 26.9020 49.9530 ;
    RECT 26.4160 49.9530 26.9020 50.0850 ;
    RECT 26.4160 50.0850 26.9020 50.1550 ;
    RECT 26.4160 50.1550 26.9660 50.7410 ;
    RECT 26.4160 50.7410 26.9020 50.8430 ;
    RECT 26.4160 50.8430 26.9020 50.9130 ;
    RECT 26.4160 50.9130 26.9020 51.0450 ;
    RECT 26.4160 51.0450 26.9020 51.1150 ;
    RECT 26.4160 51.1150 26.9660 51.7010 ;
    RECT 26.4160 51.7010 26.9020 51.8030 ;
    RECT 26.4160 51.8030 26.9020 51.8730 ;
    RECT 26.4160 51.8730 26.9020 52.0050 ;
    RECT 26.4160 52.0050 26.9020 52.0750 ;
    RECT 26.4160 52.0750 26.9660 52.6610 ;
    RECT 26.4160 52.6610 26.9020 52.7630 ;
    RECT 26.4160 52.7630 26.9020 52.8330 ;
    RECT 26.4160 52.8330 26.9020 52.9650 ;
    RECT 26.4160 52.9650 26.9020 53.0350 ;
    RECT 26.4160 53.0350 26.9660 53.6210 ;
    RECT 26.4160 53.6210 26.9020 53.7230 ;
    RECT 26.4160 53.7230 26.9020 53.7930 ;
    RECT 26.4160 53.7930 26.9020 53.9250 ;
    RECT 26.4160 53.9250 26.9020 53.9950 ;
    RECT 26.4160 53.9950 26.9660 54.5810 ;
    RECT 26.4160 54.5810 26.9020 54.6830 ;
    RECT 26.4160 54.6830 26.9020 54.7530 ;
    RECT 26.4160 54.7530 26.9020 54.8850 ;
    RECT 26.4160 54.8850 26.9020 54.9550 ;
    RECT 26.4160 54.9550 26.9660 55.5410 ;
    RECT 26.4160 55.5410 26.9020 55.6430 ;
    RECT 26.4160 55.6430 26.9020 55.7130 ;
    RECT 26.4160 55.7130 26.9020 55.8450 ;
    RECT 26.4160 55.8450 26.9020 55.9150 ;
    RECT 26.4160 55.9150 26.9660 56.5010 ;
    RECT 26.4160 56.5010 26.9020 56.6030 ;
    RECT 26.4160 56.6030 26.9020 56.6730 ;
    RECT 26.4160 56.6730 26.9020 56.8050 ;
    RECT 26.4160 56.8050 26.9020 56.8750 ;
    RECT 26.4160 56.8750 26.9660 57.4610 ;
    RECT 26.4160 57.4610 26.9020 57.5630 ;
    RECT 26.4160 57.5630 26.9020 57.6330 ;
    RECT 26.4160 57.6330 26.9020 57.7650 ;
    RECT 26.4160 57.7650 26.9020 57.8350 ;
    RECT 26.4160 57.8350 26.9660 58.4210 ;
    RECT 26.4160 58.4210 26.9020 58.5230 ;
    RECT 26.4160 58.5230 26.9020 58.5930 ;
    RECT 26.4160 58.5930 26.9020 58.7250 ;
    RECT 26.4160 58.7250 26.9020 58.7950 ;
    RECT 26.4160 58.7950 26.9660 59.3810 ;
    RECT 26.4160 59.3810 26.9020 59.4830 ;
    RECT 26.4160 59.4830 26.9020 59.5530 ;
    RECT 26.4160 59.5530 26.9020 59.6850 ;
    RECT 26.4160 59.6850 26.9020 59.7550 ;
    RECT 26.4160 59.7550 26.9660 60.3410 ;
    RECT 26.4160 60.3410 26.9020 60.4430 ;
    RECT 26.4160 60.4430 26.9020 60.5130 ;
    RECT 26.4160 60.5130 26.9020 60.6450 ;
    RECT 26.4160 60.6450 26.9020 60.7150 ;
    RECT 26.4160 60.7150 26.9660 61.3010 ;
    RECT 26.4160 61.3010 26.9020 61.4030 ;
    RECT 26.4160 61.4030 26.9020 61.4730 ;
    RECT 26.4160 61.4730 26.9020 61.6050 ;
    RECT 26.4160 61.6050 26.9020 61.6750 ;
    RECT 26.4160 61.6750 26.9660 62.2610 ;
    RECT 26.4160 62.2610 26.9020 62.3630 ;
    RECT 26.4160 62.3630 26.9020 62.4330 ;
    RECT 26.4160 62.4330 26.9020 62.5650 ;
    RECT 26.4160 62.5650 26.9020 62.6350 ;
    RECT 26.4160 62.6350 26.9660 63.2210 ;
    RECT 26.4160 63.2210 26.9020 63.3230 ;
    RECT 26.4160 63.3230 26.9020 63.3930 ;
    RECT 26.4160 63.3930 26.9020 63.5250 ;
    RECT 26.4160 63.5250 26.9020 63.5950 ;
    RECT 26.4160 63.5950 26.9660 64.1810 ;
    RECT 26.4160 64.1810 26.9020 64.2830 ;
    RECT 26.4160 64.2830 26.9020 64.3530 ;
    RECT 26.4160 64.3530 26.9020 64.4850 ;
    RECT 26.4160 64.4850 26.9020 64.5550 ;
    RECT 26.4160 64.5550 26.9660 65.1410 ;
    RECT 26.4160 65.1410 26.9020 65.2430 ;
    RECT 26.4160 65.2430 26.9020 65.3130 ;
    RECT 26.4160 65.3130 26.9020 65.4450 ;
    RECT 26.4160 65.4450 26.9020 65.5150 ;
    RECT 26.4160 65.5150 26.9660 66.1010 ;
    RECT 26.4160 66.1010 26.9020 66.2030 ;
    RECT 26.4160 66.2030 26.9020 66.2730 ;
    RECT 26.4160 66.2730 26.9020 66.4050 ;
    RECT 26.4160 66.4050 26.9020 66.4750 ;
    RECT 26.4160 66.4750 26.9660 67.0610 ;
    RECT 26.4160 67.0610 26.9020 67.1630 ;
    RECT 26.4160 67.1630 26.9020 67.2330 ;
    RECT 26.4160 67.2330 26.9020 67.3650 ;
    RECT 26.4160 67.3650 26.9020 67.4350 ;
    RECT 26.4160 67.4350 26.9660 68.0210 ;
    RECT 26.4160 68.0210 26.9020 68.1230 ;
    RECT 26.4160 68.1230 26.9020 68.1930 ;
    RECT 26.4160 68.1930 26.9020 68.3250 ;
    RECT 26.4160 68.3250 26.9020 68.3950 ;
    RECT 26.4160 68.3950 26.9660 68.9810 ;
    RECT 26.4160 68.9810 26.9020 69.0830 ;
    RECT 26.4160 69.0830 26.9020 69.1530 ;
    RECT 26.4160 69.1530 26.9020 69.2850 ;
    RECT 26.4160 69.2850 26.9020 69.3550 ;
    RECT 26.4160 69.3550 26.9660 69.9410 ;
    RECT 26.4160 69.9410 26.9020 70.0430 ;
    RECT 26.4160 70.0430 26.9020 70.1130 ;
    RECT 26.4160 70.1130 26.9020 70.2450 ;
    RECT 26.4160 70.2450 26.9020 70.3150 ;
    RECT 26.4160 70.3150 26.9660 70.9010 ;
    RECT 26.4160 70.9010 26.9020 71.0030 ;
    RECT 26.4160 71.0030 26.9020 71.0730 ;
    RECT 26.4160 71.0730 26.9020 71.2050 ;
    RECT 26.4160 71.2050 26.9020 71.2750 ;
    RECT 26.4160 71.2750 26.9660 72.0960 ;
    RECT 0.0000 0.0000 0.5500 72.0960 ;
    RECT 0.0000 0.0000 26.9660 0.5500 ;
    RECT 0.0000 71.5460 26.9660 72.0960 ;
    LAYER M4 ;
    RECT 0.0000 0.8580 14.3380 0.9670 ;
    RECT 0.0000 1.0490 14.3380 1.1580 ;
    RECT 0.0000 1.3380 14.3380 1.4470 ;
    RECT 0.0000 1.8180 14.3380 1.9270 ;
    RECT 0.0000 2.0090 14.3380 2.1180 ;
    RECT 0.0000 2.2980 14.3380 2.4070 ;
    RECT 0.0000 2.7780 14.3380 2.8870 ;
    RECT 0.0000 2.9690 14.3380 3.0780 ;
    RECT 0.0000 3.2580 14.3380 3.3670 ;
    RECT 0.0000 3.7380 14.3380 3.8470 ;
    RECT 0.0000 3.9290 14.3380 4.0380 ;
    RECT 0.0000 4.2180 14.3380 4.3270 ;
    RECT 0.0000 4.6980 14.3380 4.8070 ;
    RECT 0.0000 4.8890 14.3380 4.9980 ;
    RECT 0.0000 5.1780 14.3380 5.2870 ;
    RECT 0.0000 5.6580 14.3380 5.7670 ;
    RECT 0.0000 5.8490 14.3380 5.9580 ;
    RECT 0.0000 6.1380 14.3380 6.2470 ;
    RECT 0.0000 6.6180 14.3380 6.7270 ;
    RECT 0.0000 6.8090 14.3380 6.9180 ;
    RECT 0.0000 7.0980 14.3380 7.2070 ;
    RECT 0.0000 7.5780 14.3380 7.6870 ;
    RECT 0.0000 7.7690 14.3380 7.8780 ;
    RECT 0.0000 8.0580 14.3380 8.1670 ;
    RECT 0.0000 8.5380 14.3380 8.6470 ;
    RECT 0.0000 8.7290 14.3380 8.8380 ;
    RECT 0.0000 9.0180 14.3380 9.1270 ;
    RECT 0.0000 9.4980 14.3380 9.6070 ;
    RECT 0.0000 9.6890 14.3380 9.7980 ;
    RECT 0.0000 9.9780 14.3380 10.0870 ;
    RECT 0.0000 10.4580 14.3380 10.5670 ;
    RECT 0.0000 10.6490 14.3380 10.7580 ;
    RECT 0.0000 10.9380 14.3380 11.0470 ;
    RECT 0.0000 11.4180 14.3380 11.5270 ;
    RECT 0.0000 11.6090 14.3380 11.7180 ;
    RECT 0.0000 11.8980 14.3380 12.0070 ;
    RECT 0.0000 12.3780 14.3380 12.4870 ;
    RECT 0.0000 12.5690 14.3380 12.6780 ;
    RECT 0.0000 12.8580 14.3380 12.9670 ;
    RECT 0.0000 13.3380 14.3380 13.4470 ;
    RECT 0.0000 13.5290 14.3380 13.6380 ;
    RECT 0.0000 13.8180 14.3380 13.9270 ;
    RECT 0.0000 14.2980 14.3380 14.4070 ;
    RECT 0.0000 14.4890 14.3380 14.5980 ;
    RECT 0.0000 14.7780 14.3380 14.8870 ;
    RECT 0.0000 15.2580 14.3380 15.3670 ;
    RECT 0.0000 15.4490 14.3380 15.5580 ;
    RECT 0.0000 15.7380 14.3380 15.8470 ;
    RECT 0.0000 16.2180 14.3380 16.3270 ;
    RECT 0.0000 16.4090 14.3380 16.5180 ;
    RECT 0.0000 16.6980 14.3380 16.8070 ;
    RECT 0.0000 17.1780 14.3380 17.2870 ;
    RECT 0.0000 17.3690 14.3380 17.4780 ;
    RECT 0.0000 17.6580 14.3380 17.7670 ;
    RECT 0.0000 18.1380 14.3380 18.2470 ;
    RECT 0.0000 18.3290 14.3380 18.4380 ;
    RECT 0.0000 18.6180 14.3380 18.7270 ;
    RECT 0.0000 19.0980 14.3380 19.2070 ;
    RECT 0.0000 19.2890 14.3380 19.3980 ;
    RECT 0.0000 19.5780 14.3380 19.6870 ;
    RECT 0.0000 20.0580 14.3380 20.1670 ;
    RECT 0.0000 20.2490 14.3380 20.3580 ;
    RECT 0.0000 20.5380 14.3380 20.6470 ;
    RECT 0.0000 21.0180 14.3380 21.1270 ;
    RECT 0.0000 21.2090 14.3380 21.3180 ;
    RECT 0.0000 21.4980 14.3380 21.6070 ;
    RECT 0.0000 21.9780 14.3380 22.0870 ;
    RECT 0.0000 22.1690 14.3380 22.2780 ;
    RECT 0.0000 22.4580 14.3380 22.5670 ;
    RECT 0.0000 22.9380 14.3380 23.0470 ;
    RECT 0.0000 23.1290 14.3380 23.2380 ;
    RECT 0.0000 23.4180 14.3380 23.5270 ;
    RECT 0.0000 23.8980 14.3380 24.0070 ;
    RECT 0.0000 24.0890 14.3380 24.1980 ;
    RECT 0.0000 24.3780 14.3380 24.4870 ;
    RECT 0.0000 24.8580 14.3380 24.9670 ;
    RECT 0.0000 25.0490 14.3380 25.1580 ;
    RECT 0.0000 25.3380 14.3380 25.4470 ;
    RECT 0.0000 25.8180 14.3380 25.9270 ;
    RECT 0.0000 26.0090 14.3380 26.1180 ;
    RECT 0.0000 26.2980 14.3380 26.4070 ;
    RECT 0.0000 26.7780 14.3380 26.8870 ;
    RECT 0.0000 26.9690 14.3380 27.0780 ;
    RECT 0.0000 27.2580 14.3380 27.3670 ;
    RECT 0.0000 27.7380 14.3380 27.8470 ;
    RECT 0.0000 27.9290 14.3380 28.0380 ;
    RECT 0.0000 28.2180 14.3380 28.3270 ;
    RECT 0.0000 28.6980 14.3380 28.8070 ;
    RECT 0.0000 28.8890 14.3380 28.9980 ;
    RECT 0.0000 29.1780 14.3380 29.2870 ;
    RECT 0.0000 29.6580 14.3380 29.7670 ;
    RECT 0.0000 29.8490 14.3380 29.9580 ;
    RECT 0.0000 30.1380 14.3380 30.2470 ;
    RECT 0.0000 30.6180 14.3380 30.7270 ;
    RECT 0.0000 30.8090 14.3380 30.9180 ;
    RECT 0.0000 31.0980 14.3380 31.2070 ;
    RECT 0.0000 32.4880 16.6950 32.6080 ;
    RECT 0.0000 32.6880 16.6950 32.8080 ;
    RECT 0.0000 32.8880 16.6950 33.0080 ;
    RECT 0.0000 33.0880 16.6950 33.2080 ;
    RECT 0.0000 33.2880 16.6950 33.4080 ;
    RECT 0.0000 33.4880 16.6950 33.6080 ;
    RECT 0.0000 33.8880 16.6950 34.0080 ;
    RECT 0.0000 34.0880 16.6950 34.2080 ;
    RECT 0.0000 34.2880 16.6950 34.4080 ;
    RECT 0.0000 35.0880 16.6950 35.2080 ;
    RECT 0.0000 35.2880 16.6950 35.4080 ;
    RECT 0.0000 35.4880 16.6950 35.6080 ;
    RECT 0.0000 35.6880 16.6950 35.8080 ;
    RECT 0.0000 35.8880 16.6950 36.0080 ;
    RECT 0.0000 36.0880 15.9490 36.2080 ;
    RECT 0.0000 36.2880 16.6950 36.4080 ;
    RECT 0.0000 36.8880 16.6950 37.0080 ;
    RECT 0.0000 37.0880 16.6950 37.2080 ;
    RECT 0.0000 37.2880 16.6950 37.4080 ;
    RECT 0.0000 37.6880 16.6950 37.8080 ;
    RECT 0.0000 38.0880 16.6950 38.2080 ;
    RECT 0.0000 38.4880 16.6950 38.6080 ;
    RECT 0.0000 38.6880 16.6950 38.8080 ;
    RECT 0.0000 38.8880 16.6950 39.0080 ;
    RECT 0.0000 39.0880 16.6950 39.2080 ;
    RECT 0.0000 39.2880 16.6950 39.4080 ;
    RECT 0.0000 39.4880 16.6950 39.6080 ;
    RECT 0.0000 39.6880 16.6950 39.8080 ;
    RECT 0.0000 41.1780 14.3380 41.2870 ;
    RECT 0.0000 41.3690 14.3380 41.4780 ;
    RECT 0.0000 41.6580 14.3380 41.7670 ;
    RECT 0.0000 42.1380 14.3380 42.2470 ;
    RECT 0.0000 42.3290 14.3380 42.4380 ;
    RECT 0.0000 42.6180 14.3380 42.7270 ;
    RECT 0.0000 43.0980 14.3380 43.2070 ;
    RECT 0.0000 43.2890 14.3380 43.3980 ;
    RECT 0.0000 43.5780 14.3380 43.6870 ;
    RECT 0.0000 44.0580 14.3380 44.1670 ;
    RECT 0.0000 44.2490 14.3380 44.3580 ;
    RECT 0.0000 44.5380 14.3380 44.6470 ;
    RECT 0.0000 45.0180 14.3380 45.1270 ;
    RECT 0.0000 45.2090 14.3380 45.3180 ;
    RECT 0.0000 45.4980 14.3380 45.6070 ;
    RECT 0.0000 45.9780 14.3380 46.0870 ;
    RECT 0.0000 46.1690 14.3380 46.2780 ;
    RECT 0.0000 46.4580 14.3380 46.5670 ;
    RECT 0.0000 46.9380 14.3380 47.0470 ;
    RECT 0.0000 47.1290 14.3380 47.2380 ;
    RECT 0.0000 47.4180 14.3380 47.5270 ;
    RECT 0.0000 47.8980 14.3380 48.0070 ;
    RECT 0.0000 48.0890 14.3380 48.1980 ;
    RECT 0.0000 48.3780 14.3380 48.4870 ;
    RECT 0.0000 48.8580 14.3380 48.9670 ;
    RECT 0.0000 49.0490 14.3380 49.1580 ;
    RECT 0.0000 49.3380 14.3380 49.4470 ;
    RECT 0.0000 49.8180 14.3380 49.9270 ;
    RECT 0.0000 50.0090 14.3380 50.1180 ;
    RECT 0.0000 50.2980 14.3380 50.4070 ;
    RECT 0.0000 50.7780 14.3380 50.8870 ;
    RECT 0.0000 50.9690 14.3380 51.0780 ;
    RECT 0.0000 51.2580 14.3380 51.3670 ;
    RECT 0.0000 51.7380 14.3380 51.8470 ;
    RECT 0.0000 51.9290 14.3380 52.0380 ;
    RECT 0.0000 52.2180 14.3380 52.3270 ;
    RECT 0.0000 52.6980 14.3380 52.8070 ;
    RECT 0.0000 52.8890 14.3380 52.9980 ;
    RECT 0.0000 53.1780 14.3380 53.2870 ;
    RECT 0.0000 53.6580 14.3380 53.7670 ;
    RECT 0.0000 53.8490 14.3380 53.9580 ;
    RECT 0.0000 54.1380 14.3380 54.2470 ;
    RECT 0.0000 54.6180 14.3380 54.7270 ;
    RECT 0.0000 54.8090 14.3380 54.9180 ;
    RECT 0.0000 55.0980 14.3380 55.2070 ;
    RECT 0.0000 55.5780 14.3380 55.6870 ;
    RECT 0.0000 55.7690 14.3380 55.8780 ;
    RECT 0.0000 56.0580 14.3380 56.1670 ;
    RECT 0.0000 56.5380 14.3380 56.6470 ;
    RECT 0.0000 56.7290 14.3380 56.8380 ;
    RECT 0.0000 57.0180 14.3380 57.1270 ;
    RECT 0.0000 57.4980 14.3380 57.6070 ;
    RECT 0.0000 57.6890 14.3380 57.7980 ;
    RECT 0.0000 57.9780 14.3380 58.0870 ;
    RECT 0.0000 58.4580 14.3380 58.5670 ;
    RECT 0.0000 58.6490 14.3380 58.7580 ;
    RECT 0.0000 58.9380 14.3380 59.0470 ;
    RECT 0.0000 59.4180 14.3380 59.5270 ;
    RECT 0.0000 59.6090 14.3380 59.7180 ;
    RECT 0.0000 59.8980 14.3380 60.0070 ;
    RECT 0.0000 60.3780 14.3380 60.4870 ;
    RECT 0.0000 60.5690 14.3380 60.6780 ;
    RECT 0.0000 60.8580 14.3380 60.9670 ;
    RECT 0.0000 61.3380 14.3380 61.4470 ;
    RECT 0.0000 61.5290 14.3380 61.6380 ;
    RECT 0.0000 61.8180 14.3380 61.9270 ;
    RECT 0.0000 62.2980 14.3380 62.4070 ;
    RECT 0.0000 62.4890 14.3380 62.5980 ;
    RECT 0.0000 62.7780 14.3380 62.8870 ;
    RECT 0.0000 63.2580 14.3380 63.3670 ;
    RECT 0.0000 63.4490 14.3380 63.5580 ;
    RECT 0.0000 63.7380 14.3380 63.8470 ;
    RECT 0.0000 64.2180 14.3380 64.3270 ;
    RECT 0.0000 64.4090 14.3380 64.5180 ;
    RECT 0.0000 64.6980 14.3380 64.8070 ;
    RECT 0.0000 65.1780 14.3380 65.2870 ;
    RECT 0.0000 65.3690 14.3380 65.4780 ;
    RECT 0.0000 65.6580 14.3380 65.7670 ;
    RECT 0.0000 66.1380 14.3380 66.2470 ;
    RECT 0.0000 66.3290 14.3380 66.4380 ;
    RECT 0.0000 66.6180 14.3380 66.7270 ;
    RECT 0.0000 67.0980 14.3380 67.2070 ;
    RECT 0.0000 67.2890 14.3380 67.3980 ;
    RECT 0.0000 67.5780 14.3380 67.6870 ;
    RECT 0.0000 68.0580 14.3380 68.1670 ;
    RECT 0.0000 68.2490 14.3380 68.3580 ;
    RECT 0.0000 68.5380 14.3380 68.6470 ;
    RECT 0.0000 69.0180 14.3380 69.1270 ;
    RECT 0.0000 69.2090 14.3380 69.3180 ;
    RECT 0.0000 69.4980 14.3380 69.6070 ;
    RECT 0.0000 69.9780 14.3380 70.0870 ;
    RECT 0.0000 70.1690 14.3380 70.2780 ;
    RECT 0.0000 70.4580 14.3380 70.5670 ;
    RECT 0.0000 70.9380 14.3380 71.0470 ;
    RECT 0.0000 71.1290 14.3380 71.2380 ;
    RECT 0.0000 71.4180 14.3380 71.5270 ;
  END
  PIN VDD
  USE POWER ;
  DIRECTION INOUT ;
    PORT
      LAYER M4 ;
      RECT 0.0000 0.5690 26.7280 0.6780 ;
      RECT 14.4780 1.0490 26.7280 1.1580 ;
      RECT 0.0000 1.5290 14.3380 1.6380 ;
      RECT 14.4780 1.5290 26.7280 1.6380 ;
      RECT 14.4780 2.0090 26.7280 2.1180 ;
      RECT 0.0000 2.4890 26.7280 2.5980 ;
      RECT 14.4780 2.9690 26.7280 3.0780 ;
      RECT 0.0000 3.4490 14.3380 3.5580 ;
      RECT 14.4780 3.4490 26.7280 3.5580 ;
      RECT 14.4780 3.9290 26.7280 4.0380 ;
      RECT 0.0000 4.4090 26.7280 4.5180 ;
      RECT 14.4780 4.8890 26.7280 4.9980 ;
      RECT 0.0000 5.3690 14.3380 5.4780 ;
      RECT 14.4780 5.3690 26.7280 5.4780 ;
      RECT 14.4780 5.8490 26.7280 5.9580 ;
      RECT 0.0000 6.3290 26.7280 6.4380 ;
      RECT 14.4780 6.8090 26.7280 6.9180 ;
      RECT 0.0000 7.2890 14.3380 7.3980 ;
      RECT 14.4780 7.2890 26.7280 7.3980 ;
      RECT 14.4780 7.7690 26.7280 7.8780 ;
      RECT 0.0000 8.2490 26.7280 8.3580 ;
      RECT 14.4780 8.7290 26.7280 8.8380 ;
      RECT 0.0000 9.2090 14.3380 9.3180 ;
      RECT 14.4780 9.2090 26.7280 9.3180 ;
      RECT 14.4780 9.6890 26.7280 9.7980 ;
      RECT 0.0000 10.1690 26.7280 10.2780 ;
      RECT 14.4780 10.6490 26.7280 10.7580 ;
      RECT 0.0000 11.1290 14.3380 11.2380 ;
      RECT 14.4780 11.1290 26.7280 11.2380 ;
      RECT 14.4780 11.6090 26.7280 11.7180 ;
      RECT 0.0000 12.0890 26.7280 12.1980 ;
      RECT 14.4780 12.5690 26.7280 12.6780 ;
      RECT 0.0000 13.0490 14.3380 13.1580 ;
      RECT 14.4780 13.0490 26.7280 13.1580 ;
      RECT 14.4780 13.5290 26.7280 13.6380 ;
      RECT 0.0000 14.0090 26.7280 14.1180 ;
      RECT 14.4780 14.4890 26.7280 14.5980 ;
      RECT 0.0000 14.9690 14.3380 15.0780 ;
      RECT 14.4780 14.9690 26.7280 15.0780 ;
      RECT 14.4780 15.4490 26.7280 15.5580 ;
      RECT 0.0000 15.9290 26.7280 16.0380 ;
      RECT 14.4780 16.4090 26.7280 16.5180 ;
      RECT 0.0000 16.8890 14.3380 16.9980 ;
      RECT 14.4780 16.8890 26.7280 16.9980 ;
      RECT 14.4780 17.3690 26.7280 17.4780 ;
      RECT 0.0000 17.8490 26.7280 17.9580 ;
      RECT 14.4780 18.3290 26.7280 18.4380 ;
      RECT 0.0000 18.8090 14.3380 18.9180 ;
      RECT 14.4780 18.8090 26.7280 18.9180 ;
      RECT 14.4780 19.2890 26.7280 19.3980 ;
      RECT 0.0000 19.7690 26.7280 19.8780 ;
      RECT 14.4780 20.2490 26.7280 20.3580 ;
      RECT 0.0000 20.7290 14.3380 20.8380 ;
      RECT 14.4780 20.7290 26.7280 20.8380 ;
      RECT 14.4780 21.2090 26.7280 21.3180 ;
      RECT 0.0000 21.6890 26.7280 21.7980 ;
      RECT 14.4780 22.1690 26.7280 22.2780 ;
      RECT 0.0000 22.6490 14.3380 22.7580 ;
      RECT 14.4780 22.6490 26.7280 22.7580 ;
      RECT 14.4780 23.1290 26.7280 23.2380 ;
      RECT 0.0000 23.6090 26.7280 23.7180 ;
      RECT 14.4780 24.0890 26.7280 24.1980 ;
      RECT 0.0000 24.5690 14.3380 24.6780 ;
      RECT 14.4780 24.5690 26.7280 24.6780 ;
      RECT 14.4780 25.0490 26.7280 25.1580 ;
      RECT 0.0000 25.5290 26.7280 25.6380 ;
      RECT 14.4780 26.0090 26.7280 26.1180 ;
      RECT 0.0000 26.4890 14.3380 26.5980 ;
      RECT 14.4780 26.4890 26.7280 26.5980 ;
      RECT 14.4780 26.9690 26.7280 27.0780 ;
      RECT 0.0000 27.4490 26.7280 27.5580 ;
      RECT 14.4780 27.9290 26.7280 28.0380 ;
      RECT 0.0000 28.4090 14.3380 28.5180 ;
      RECT 14.4780 28.4090 26.7280 28.5180 ;
      RECT 14.4780 28.8890 26.7280 28.9980 ;
      RECT 0.0000 29.3690 26.7280 29.4780 ;
      RECT 14.4780 29.8490 26.7280 29.9580 ;
      RECT 0.0000 30.3290 14.3380 30.4380 ;
      RECT 14.4780 30.3290 26.7280 30.4380 ;
      RECT 14.4780 30.8090 26.7280 30.9180 ;
      RECT 16.8350 32.4880 26.7520 32.6080 ;
      RECT 16.8350 32.6880 26.7520 32.8080 ;
      RECT 16.8350 32.8880 26.7520 33.0080 ;
      RECT 16.8350 33.0880 26.7520 33.2080 ;
      RECT 16.8350 33.2880 26.7520 33.4080 ;
      RECT 16.8350 33.4880 26.7520 33.6080 ;
      RECT 0.0000 33.6880 16.6950 33.8080 ;
      RECT 16.8350 33.6880 26.7520 33.8080 ;
      RECT 16.8350 33.8880 26.7520 34.0080 ;
      RECT 16.8350 34.2880 26.7520 34.4080 ;
      RECT 0.0000 34.4880 16.6950 34.6080 ;
      RECT 16.8350 34.6880 26.7520 34.8080 ;
      RECT 16.8350 35.0880 26.7520 35.2080 ;
      RECT 16.8350 35.4880 26.7520 35.6080 ;
      RECT 16.8350 35.8880 26.7520 36.0080 ;
      RECT 16.8350 36.2880 26.7520 36.4080 ;
      RECT 16.8350 36.6880 26.7520 36.8080 ;
      RECT 16.8350 37.0880 26.7520 37.2080 ;
      RECT 0.0000 37.4880 16.6950 37.6080 ;
      RECT 16.8350 37.4880 26.7520 37.6080 ;
      RECT 16.8350 37.8880 26.7520 38.0080 ;
      RECT 0.0000 38.2880 16.6950 38.4080 ;
      RECT 16.8350 38.2880 26.7520 38.4080 ;
      RECT 16.8350 38.6880 26.7520 38.8080 ;
      RECT 16.8350 38.8880 26.7520 39.0080 ;
      RECT 16.8350 39.0880 26.7520 39.2080 ;
      RECT 16.8350 39.2880 26.7520 39.4080 ;
      RECT 16.8350 39.4880 26.7520 39.6080 ;
      RECT 0.0000 40.8890 26.7280 40.9980 ;
      RECT 14.4780 41.3690 26.7280 41.4780 ;
      RECT 0.0000 41.8490 14.3380 41.9580 ;
      RECT 14.4780 41.8490 26.7280 41.9580 ;
      RECT 14.4780 42.3290 26.7280 42.4380 ;
      RECT 0.0000 42.8090 26.7280 42.9180 ;
      RECT 14.4780 43.2890 26.7280 43.3980 ;
      RECT 0.0000 43.7690 14.3380 43.8780 ;
      RECT 14.4780 43.7690 26.7280 43.8780 ;
      RECT 14.4780 44.2490 26.7280 44.3580 ;
      RECT 0.0000 44.7290 26.7280 44.8380 ;
      RECT 14.4780 45.2090 26.7280 45.3180 ;
      RECT 0.0000 45.6890 14.3380 45.7980 ;
      RECT 14.4780 45.6890 26.7280 45.7980 ;
      RECT 14.4780 46.1690 26.7280 46.2780 ;
      RECT 0.0000 46.6490 26.7280 46.7580 ;
      RECT 14.4780 47.1290 26.7280 47.2380 ;
      RECT 0.0000 47.6090 14.3380 47.7180 ;
      RECT 14.4780 47.6090 26.7280 47.7180 ;
      RECT 14.4780 48.0890 26.7280 48.1980 ;
      RECT 0.0000 48.5690 26.7280 48.6780 ;
      RECT 14.4780 49.0490 26.7280 49.1580 ;
      RECT 0.0000 49.5290 14.3380 49.6380 ;
      RECT 14.4780 49.5290 26.7280 49.6380 ;
      RECT 14.4780 50.0090 26.7280 50.1180 ;
      RECT 0.0000 50.4890 26.7280 50.5980 ;
      RECT 14.4780 50.9690 26.7280 51.0780 ;
      RECT 0.0000 51.4490 14.3380 51.5580 ;
      RECT 14.4780 51.4490 26.7280 51.5580 ;
      RECT 14.4780 51.9290 26.7280 52.0380 ;
      RECT 0.0000 52.4090 26.7280 52.5180 ;
      RECT 14.4780 52.8890 26.7280 52.9980 ;
      RECT 0.0000 53.3690 14.3380 53.4780 ;
      RECT 14.4780 53.3690 26.7280 53.4780 ;
      RECT 14.4780 53.8490 26.7280 53.9580 ;
      RECT 0.0000 54.3290 26.7280 54.4380 ;
      RECT 14.4780 54.8090 26.7280 54.9180 ;
      RECT 0.0000 55.2890 14.3380 55.3980 ;
      RECT 14.4780 55.2890 26.7280 55.3980 ;
      RECT 14.4780 55.7690 26.7280 55.8780 ;
      RECT 0.0000 56.2490 26.7280 56.3580 ;
      RECT 14.4780 56.7290 26.7280 56.8380 ;
      RECT 0.0000 57.2090 14.3380 57.3180 ;
      RECT 14.4780 57.2090 26.7280 57.3180 ;
      RECT 14.4780 57.6890 26.7280 57.7980 ;
      RECT 0.0000 58.1690 26.7280 58.2780 ;
      RECT 14.4780 58.6490 26.7280 58.7580 ;
      RECT 0.0000 59.1290 14.3380 59.2380 ;
      RECT 14.4780 59.1290 26.7280 59.2380 ;
      RECT 14.4780 59.6090 26.7280 59.7180 ;
      RECT 0.0000 60.0890 26.7280 60.1980 ;
      RECT 14.4780 60.5690 26.7280 60.6780 ;
      RECT 0.0000 61.0490 14.3380 61.1580 ;
      RECT 14.4780 61.0490 26.7280 61.1580 ;
      RECT 14.4780 61.5290 26.7280 61.6380 ;
      RECT 0.0000 62.0090 26.7280 62.1180 ;
      RECT 14.4780 62.4890 26.7280 62.5980 ;
      RECT 0.0000 62.9690 14.3380 63.0780 ;
      RECT 14.4780 62.9690 26.7280 63.0780 ;
      RECT 14.4780 63.4490 26.7280 63.5580 ;
      RECT 0.0000 63.9290 26.7280 64.0380 ;
      RECT 14.4780 64.4090 26.7280 64.5180 ;
      RECT 0.0000 64.8890 14.3380 64.9980 ;
      RECT 14.4780 64.8890 26.7280 64.9980 ;
      RECT 14.4780 65.3690 26.7280 65.4780 ;
      RECT 0.0000 65.8490 26.7280 65.9580 ;
      RECT 14.4780 66.3290 26.7280 66.4380 ;
      RECT 0.0000 66.8090 14.3380 66.9180 ;
      RECT 14.4780 66.8090 26.7280 66.9180 ;
      RECT 14.4780 67.2890 26.7280 67.3980 ;
      RECT 0.0000 67.7690 26.7280 67.8780 ;
      RECT 14.4780 68.2490 26.7280 68.3580 ;
      RECT 0.0000 68.7290 14.3380 68.8380 ;
      RECT 14.4780 68.7290 26.7280 68.8380 ;
      RECT 14.4780 69.2090 26.7280 69.3180 ;
      RECT 0.0000 69.6890 26.7280 69.7980 ;
      RECT 14.4780 70.1690 26.7280 70.2780 ;
      RECT 0.0000 70.6490 14.3380 70.7580 ;
      RECT 14.4780 70.6490 26.7280 70.7580 ;
      RECT 14.4780 71.1290 26.7280 71.2380 ;
    END
  END VDD
  PIN VSS
  USE GROUND ;
  DIRECTION INOUT ;
    PORT
      LAYER M4 ;
      RECT 14.4780 0.8580 26.7280 0.9670 ;
      RECT 14.4780 1.3380 26.7280 1.4470 ;
      RECT 14.4780 1.8180 26.7280 1.9270 ;
      RECT 14.4780 2.2980 26.7280 2.4070 ;
      RECT 14.4780 2.7780 26.7280 2.8870 ;
      RECT 14.4780 3.2580 26.7280 3.3670 ;
      RECT 14.4780 3.7380 26.7280 3.8470 ;
      RECT 14.4780 4.2180 26.7280 4.3270 ;
      RECT 14.4780 4.6980 26.7280 4.8070 ;
      RECT 14.4780 5.1780 26.7280 5.2870 ;
      RECT 14.4780 5.6580 26.7280 5.7670 ;
      RECT 14.4780 6.1380 26.7280 6.2470 ;
      RECT 14.4780 6.6180 26.7280 6.7270 ;
      RECT 14.4780 7.0980 26.7280 7.2070 ;
      RECT 14.4780 7.5780 26.7280 7.6870 ;
      RECT 14.4780 8.0580 26.7280 8.1670 ;
      RECT 14.4780 8.5380 26.7280 8.6470 ;
      RECT 14.4780 9.0180 26.7280 9.1270 ;
      RECT 14.4780 9.4980 26.7280 9.6070 ;
      RECT 14.4780 9.9780 26.7280 10.0870 ;
      RECT 14.4780 10.4580 26.7280 10.5670 ;
      RECT 14.4780 10.9380 26.7280 11.0470 ;
      RECT 14.4780 11.4180 26.7280 11.5270 ;
      RECT 14.4780 11.8980 26.7280 12.0070 ;
      RECT 14.4780 12.3780 26.7280 12.4870 ;
      RECT 14.4780 12.8580 26.7280 12.9670 ;
      RECT 14.4780 13.3380 26.7280 13.4470 ;
      RECT 14.4780 13.8180 26.7280 13.9270 ;
      RECT 14.4780 14.2980 26.7280 14.4070 ;
      RECT 14.4780 14.7780 26.7280 14.8870 ;
      RECT 14.4780 15.2580 26.7280 15.3670 ;
      RECT 14.4780 15.7380 26.7280 15.8470 ;
      RECT 14.4780 16.2180 26.7280 16.3270 ;
      RECT 14.4780 16.6980 26.7280 16.8070 ;
      RECT 14.4780 17.1780 26.7280 17.2870 ;
      RECT 14.4780 17.6580 26.7280 17.7670 ;
      RECT 14.4780 18.1380 26.7280 18.2470 ;
      RECT 14.4780 18.6180 26.7280 18.7270 ;
      RECT 14.4780 19.0980 26.7280 19.2070 ;
      RECT 14.4780 19.5780 26.7280 19.6870 ;
      RECT 14.4780 20.0580 26.7280 20.1670 ;
      RECT 14.4780 20.5380 26.7280 20.6470 ;
      RECT 14.4780 21.0180 26.7280 21.1270 ;
      RECT 14.4780 21.4980 26.7280 21.6070 ;
      RECT 14.4780 21.9780 26.7280 22.0870 ;
      RECT 14.4780 22.4580 26.7280 22.5670 ;
      RECT 14.4780 22.9380 26.7280 23.0470 ;
      RECT 14.4780 23.4180 26.7280 23.5270 ;
      RECT 14.4780 23.8980 26.7280 24.0070 ;
      RECT 14.4780 24.3780 26.7280 24.4870 ;
      RECT 14.4780 24.8580 26.7280 24.9670 ;
      RECT 14.4780 25.3380 26.7280 25.4470 ;
      RECT 14.4780 25.8180 26.7280 25.9270 ;
      RECT 14.4780 26.2980 26.7280 26.4070 ;
      RECT 14.4780 26.7780 26.7280 26.8870 ;
      RECT 14.4780 27.2580 26.7280 27.3670 ;
      RECT 14.4780 27.7380 26.7280 27.8470 ;
      RECT 14.4780 28.2180 26.7280 28.3270 ;
      RECT 14.4780 28.6980 26.7280 28.8070 ;
      RECT 14.4780 29.1780 26.7280 29.2870 ;
      RECT 14.4780 29.6580 26.7280 29.7670 ;
      RECT 14.4780 30.1380 26.7280 30.2470 ;
      RECT 14.4780 30.6180 26.7280 30.7270 ;
      RECT 14.4780 31.0980 26.7280 31.2070 ;
      RECT 0.0000 31.2890 26.7520 31.4010 ;
      RECT 0.0000 31.6880 26.7520 31.8080 ;
      RECT 0.0000 31.8880 26.7520 32.0080 ;
      RECT 0.0000 32.0880 26.7520 32.2080 ;
      RECT 0.0000 32.2880 16.6950 32.4080 ;
      RECT 16.8350 32.2880 26.7520 32.4080 ;
      RECT 16.8350 34.0880 26.7520 34.2080 ;
      RECT 16.8350 34.4880 26.7520 34.6080 ;
      RECT 0.0000 34.6880 16.6950 34.8080 ;
      RECT 0.0000 34.8880 26.7520 35.0080 ;
      RECT 16.8350 35.2880 26.7520 35.4080 ;
      RECT 16.8350 35.6880 26.7520 35.8080 ;
      RECT 16.0890 36.0880 26.7520 36.2080 ;
      RECT 0.0000 36.4880 26.7520 36.6080 ;
      RECT 0.0000 36.6880 16.6950 36.8080 ;
      RECT 16.8350 36.8880 26.7520 37.0080 ;
      RECT 16.8350 37.2880 26.7520 37.4080 ;
      RECT 16.8350 37.6880 26.7520 37.8080 ;
      RECT 0.0000 37.8880 16.6950 38.0080 ;
      RECT 16.8350 38.0880 26.7520 38.2080 ;
      RECT 16.8350 38.4880 26.7520 38.6080 ;
      RECT 16.8350 39.6880 26.7520 39.8080 ;
      RECT 0.0000 39.8880 26.7520 40.0080 ;
      RECT 0.0000 40.0880 16.6950 40.2080 ;
      RECT 16.8350 40.0880 26.7520 40.2080 ;
      RECT 0.0000 40.2880 26.7520 40.4080 ;
      RECT 0.0000 40.6950 26.7520 40.8070 ;
      RECT 14.4780 41.1780 26.7280 41.2870 ;
      RECT 14.4780 41.6580 26.7280 41.7670 ;
      RECT 14.4780 42.1380 26.7280 42.2470 ;
      RECT 14.4780 42.6180 26.7280 42.7270 ;
      RECT 14.4780 43.0980 26.7280 43.2070 ;
      RECT 14.4780 43.5780 26.7280 43.6870 ;
      RECT 14.4780 44.0580 26.7280 44.1670 ;
      RECT 14.4780 44.5380 26.7280 44.6470 ;
      RECT 14.4780 45.0180 26.7280 45.1270 ;
      RECT 14.4780 45.4980 26.7280 45.6070 ;
      RECT 14.4780 45.9780 26.7280 46.0870 ;
      RECT 14.4780 46.4580 26.7280 46.5670 ;
      RECT 14.4780 46.9380 26.7280 47.0470 ;
      RECT 14.4780 47.4180 26.7280 47.5270 ;
      RECT 14.4780 47.8980 26.7280 48.0070 ;
      RECT 14.4780 48.3780 26.7280 48.4870 ;
      RECT 14.4780 48.8580 26.7280 48.9670 ;
      RECT 14.4780 49.3380 26.7280 49.4470 ;
      RECT 14.4780 49.8180 26.7280 49.9270 ;
      RECT 14.4780 50.2980 26.7280 50.4070 ;
      RECT 14.4780 50.7780 26.7280 50.8870 ;
      RECT 14.4780 51.2580 26.7280 51.3670 ;
      RECT 14.4780 51.7380 26.7280 51.8470 ;
      RECT 14.4780 52.2180 26.7280 52.3270 ;
      RECT 14.4780 52.6980 26.7280 52.8070 ;
      RECT 14.4780 53.1780 26.7280 53.2870 ;
      RECT 14.4780 53.6580 26.7280 53.7670 ;
      RECT 14.4780 54.1380 26.7280 54.2470 ;
      RECT 14.4780 54.6180 26.7280 54.7270 ;
      RECT 14.4780 55.0980 26.7280 55.2070 ;
      RECT 14.4780 55.5780 26.7280 55.6870 ;
      RECT 14.4780 56.0580 26.7280 56.1670 ;
      RECT 14.4780 56.5380 26.7280 56.6470 ;
      RECT 14.4780 57.0180 26.7280 57.1270 ;
      RECT 14.4780 57.4980 26.7280 57.6070 ;
      RECT 14.4780 57.9780 26.7280 58.0870 ;
      RECT 14.4780 58.4580 26.7280 58.5670 ;
      RECT 14.4780 58.9380 26.7280 59.0470 ;
      RECT 14.4780 59.4180 26.7280 59.5270 ;
      RECT 14.4780 59.8980 26.7280 60.0070 ;
      RECT 14.4780 60.3780 26.7280 60.4870 ;
      RECT 14.4780 60.8580 26.7280 60.9670 ;
      RECT 14.4780 61.3380 26.7280 61.4470 ;
      RECT 14.4780 61.8180 26.7280 61.9270 ;
      RECT 14.4780 62.2980 26.7280 62.4070 ;
      RECT 14.4780 62.7780 26.7280 62.8870 ;
      RECT 14.4780 63.2580 26.7280 63.3670 ;
      RECT 14.4780 63.7380 26.7280 63.8470 ;
      RECT 14.4780 64.2180 26.7280 64.3270 ;
      RECT 14.4780 64.6980 26.7280 64.8070 ;
      RECT 14.4780 65.1780 26.7280 65.2870 ;
      RECT 14.4780 65.6580 26.7280 65.7670 ;
      RECT 14.4780 66.1380 26.7280 66.2470 ;
      RECT 14.4780 66.6180 26.7280 66.7270 ;
      RECT 14.4780 67.0980 26.7280 67.2070 ;
      RECT 14.4780 67.5780 26.7280 67.6870 ;
      RECT 14.4780 68.0580 26.7280 68.1670 ;
      RECT 14.4780 68.5380 26.7280 68.6470 ;
      RECT 14.4780 69.0180 26.7280 69.1270 ;
      RECT 14.4780 69.4980 26.7280 69.6070 ;
      RECT 14.4780 69.9780 26.7280 70.0870 ;
      RECT 14.4780 70.4580 26.7280 70.5670 ;
      RECT 14.4780 70.9380 26.7280 71.0470 ;
      RECT 14.4780 71.4180 26.7280 71.5270 ;
    END
  END VSS
  END dti_1pr_ll_tm16ffcllhvt_64x128_1ww2x_m_shc
END LIBRARY
